// adaptor2x2.v

// Generated using ACDS version 17.1 590

`timescale 1 ps / 1 ps
module adaptor2x2 (
		input  wire  clk_clk,       //   clk.clk
		input  wire  reset_reset_n  // reset.reset_n
	);

	wire  [31:0] nios2_gen2_00_data_master_readdata;                           // mm_interconnect_0:nios2_gen2_00_data_master_readdata -> nios2_gen2_00:d_readdata
	wire         nios2_gen2_00_data_master_waitrequest;                        // mm_interconnect_0:nios2_gen2_00_data_master_waitrequest -> nios2_gen2_00:d_waitrequest
	wire         nios2_gen2_00_data_master_debugaccess;                        // nios2_gen2_00:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_00_data_master_debugaccess
	wire  [13:0] nios2_gen2_00_data_master_address;                            // nios2_gen2_00:d_address -> mm_interconnect_0:nios2_gen2_00_data_master_address
	wire   [3:0] nios2_gen2_00_data_master_byteenable;                         // nios2_gen2_00:d_byteenable -> mm_interconnect_0:nios2_gen2_00_data_master_byteenable
	wire         nios2_gen2_00_data_master_read;                               // nios2_gen2_00:d_read -> mm_interconnect_0:nios2_gen2_00_data_master_read
	wire         nios2_gen2_00_data_master_write;                              // nios2_gen2_00:d_write -> mm_interconnect_0:nios2_gen2_00_data_master_write
	wire  [31:0] nios2_gen2_00_data_master_writedata;                          // nios2_gen2_00:d_writedata -> mm_interconnect_0:nios2_gen2_00_data_master_writedata
	wire  [31:0] nios2_gen2_00_instruction_master_readdata;                    // mm_interconnect_0:nios2_gen2_00_instruction_master_readdata -> nios2_gen2_00:i_readdata
	wire         nios2_gen2_00_instruction_master_waitrequest;                 // mm_interconnect_0:nios2_gen2_00_instruction_master_waitrequest -> nios2_gen2_00:i_waitrequest
	wire  [13:0] nios2_gen2_00_instruction_master_address;                     // nios2_gen2_00:i_address -> mm_interconnect_0:nios2_gen2_00_instruction_master_address
	wire         nios2_gen2_00_instruction_master_read;                        // nios2_gen2_00:i_read -> mm_interconnect_0:nios2_gen2_00_instruction_master_read
	wire   [7:0] mm_interconnect_0_adaptor_2x2_0_input_00_readdata;            // adaptor_2x2_0:reaData_00 -> mm_interconnect_0:adaptor_2x2_0_Input_00_readdata
	wire         mm_interconnect_0_adaptor_2x2_0_input_00_read;                // mm_interconnect_0:adaptor_2x2_0_Input_00_read -> adaptor_2x2_0:read_00
	wire         mm_interconnect_0_adaptor_2x2_0_output_00_waitrequest;        // adaptor_2x2_0:waiteRequest_00 -> mm_interconnect_0:adaptor_2x2_0_Output_00_waitrequest
	wire         mm_interconnect_0_adaptor_2x2_0_output_00_write;              // mm_interconnect_0:adaptor_2x2_0_Output_00_write -> adaptor_2x2_0:write_00
	wire   [7:0] mm_interconnect_0_adaptor_2x2_0_output_00_writedata;          // mm_interconnect_0:adaptor_2x2_0_Output_00_writedata -> adaptor_2x2_0:writeData_00
	wire         mm_interconnect_0_jtag_uart_00_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_00_avalon_jtag_slave_chipselect -> jtag_uart_00:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_00_avalon_jtag_slave_readdata;    // jtag_uart_00:av_readdata -> mm_interconnect_0:jtag_uart_00_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_00_avalon_jtag_slave_waitrequest; // jtag_uart_00:av_waitrequest -> mm_interconnect_0:jtag_uart_00_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_00_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_00_avalon_jtag_slave_address -> jtag_uart_00:av_address
	wire         mm_interconnect_0_jtag_uart_00_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_00_avalon_jtag_slave_read -> jtag_uart_00:av_read_n
	wire         mm_interconnect_0_jtag_uart_00_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_00_avalon_jtag_slave_write -> jtag_uart_00:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_00_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_00_avalon_jtag_slave_writedata -> jtag_uart_00:av_writedata
	wire  [31:0] mm_interconnect_0_nios2_gen2_00_debug_mem_slave_readdata;     // nios2_gen2_00:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_00_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_00_debug_mem_slave_waitrequest;  // nios2_gen2_00:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_00_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_00_debug_mem_slave_debugaccess;  // mm_interconnect_0:nios2_gen2_00_debug_mem_slave_debugaccess -> nios2_gen2_00:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_00_debug_mem_slave_address;      // mm_interconnect_0:nios2_gen2_00_debug_mem_slave_address -> nios2_gen2_00:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_00_debug_mem_slave_read;         // mm_interconnect_0:nios2_gen2_00_debug_mem_slave_read -> nios2_gen2_00:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_00_debug_mem_slave_byteenable;   // mm_interconnect_0:nios2_gen2_00_debug_mem_slave_byteenable -> nios2_gen2_00:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_00_debug_mem_slave_write;        // mm_interconnect_0:nios2_gen2_00_debug_mem_slave_write -> nios2_gen2_00:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_00_debug_mem_slave_writedata;    // mm_interconnect_0:nios2_gen2_00_debug_mem_slave_writedata -> nios2_gen2_00:debug_mem_slave_writedata
	wire         mm_interconnect_0_data_memory_00_s1_chipselect;               // mm_interconnect_0:Data_Memory_00_s1_chipselect -> Data_Memory_00:chipselect
	wire  [31:0] mm_interconnect_0_data_memory_00_s1_readdata;                 // Data_Memory_00:readdata -> mm_interconnect_0:Data_Memory_00_s1_readdata
	wire   [9:0] mm_interconnect_0_data_memory_00_s1_address;                  // mm_interconnect_0:Data_Memory_00_s1_address -> Data_Memory_00:address
	wire   [3:0] mm_interconnect_0_data_memory_00_s1_byteenable;               // mm_interconnect_0:Data_Memory_00_s1_byteenable -> Data_Memory_00:byteenable
	wire         mm_interconnect_0_data_memory_00_s1_write;                    // mm_interconnect_0:Data_Memory_00_s1_write -> Data_Memory_00:write
	wire  [31:0] mm_interconnect_0_data_memory_00_s1_writedata;                // mm_interconnect_0:Data_Memory_00_s1_writedata -> Data_Memory_00:writedata
	wire         mm_interconnect_0_data_memory_00_s1_clken;                    // mm_interconnect_0:Data_Memory_00_s1_clken -> Data_Memory_00:clken
	wire         mm_interconnect_0_instruction_memory_00_s1_chipselect;        // mm_interconnect_0:Instruction_Memory_00_s1_chipselect -> Instruction_Memory_00:chipselect
	wire  [31:0] mm_interconnect_0_instruction_memory_00_s1_readdata;          // Instruction_Memory_00:readdata -> mm_interconnect_0:Instruction_Memory_00_s1_readdata
	wire   [9:0] mm_interconnect_0_instruction_memory_00_s1_address;           // mm_interconnect_0:Instruction_Memory_00_s1_address -> Instruction_Memory_00:address
	wire   [3:0] mm_interconnect_0_instruction_memory_00_s1_byteenable;        // mm_interconnect_0:Instruction_Memory_00_s1_byteenable -> Instruction_Memory_00:byteenable
	wire         mm_interconnect_0_instruction_memory_00_s1_write;             // mm_interconnect_0:Instruction_Memory_00_s1_write -> Instruction_Memory_00:write
	wire  [31:0] mm_interconnect_0_instruction_memory_00_s1_writedata;         // mm_interconnect_0:Instruction_Memory_00_s1_writedata -> Instruction_Memory_00:writedata
	wire         mm_interconnect_0_instruction_memory_00_s1_clken;             // mm_interconnect_0:Instruction_Memory_00_s1_clken -> Instruction_Memory_00:clken
	wire  [31:0] nios2_gen2_01_data_master_readdata;                           // mm_interconnect_1:nios2_gen2_01_data_master_readdata -> nios2_gen2_01:d_readdata
	wire         nios2_gen2_01_data_master_waitrequest;                        // mm_interconnect_1:nios2_gen2_01_data_master_waitrequest -> nios2_gen2_01:d_waitrequest
	wire         nios2_gen2_01_data_master_debugaccess;                        // nios2_gen2_01:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_1:nios2_gen2_01_data_master_debugaccess
	wire  [13:0] nios2_gen2_01_data_master_address;                            // nios2_gen2_01:d_address -> mm_interconnect_1:nios2_gen2_01_data_master_address
	wire   [3:0] nios2_gen2_01_data_master_byteenable;                         // nios2_gen2_01:d_byteenable -> mm_interconnect_1:nios2_gen2_01_data_master_byteenable
	wire         nios2_gen2_01_data_master_read;                               // nios2_gen2_01:d_read -> mm_interconnect_1:nios2_gen2_01_data_master_read
	wire         nios2_gen2_01_data_master_write;                              // nios2_gen2_01:d_write -> mm_interconnect_1:nios2_gen2_01_data_master_write
	wire  [31:0] nios2_gen2_01_data_master_writedata;                          // nios2_gen2_01:d_writedata -> mm_interconnect_1:nios2_gen2_01_data_master_writedata
	wire  [31:0] nios2_gen2_01_instruction_master_readdata;                    // mm_interconnect_1:nios2_gen2_01_instruction_master_readdata -> nios2_gen2_01:i_readdata
	wire         nios2_gen2_01_instruction_master_waitrequest;                 // mm_interconnect_1:nios2_gen2_01_instruction_master_waitrequest -> nios2_gen2_01:i_waitrequest
	wire  [13:0] nios2_gen2_01_instruction_master_address;                     // nios2_gen2_01:i_address -> mm_interconnect_1:nios2_gen2_01_instruction_master_address
	wire         nios2_gen2_01_instruction_master_read;                        // nios2_gen2_01:i_read -> mm_interconnect_1:nios2_gen2_01_instruction_master_read
	wire   [7:0] mm_interconnect_1_adaptor_2x2_0_input_01_readdata;            // adaptor_2x2_0:reaData_01 -> mm_interconnect_1:adaptor_2x2_0_Input_01_readdata
	wire         mm_interconnect_1_adaptor_2x2_0_input_01_read;                // mm_interconnect_1:adaptor_2x2_0_Input_01_read -> adaptor_2x2_0:read_01
	wire         mm_interconnect_1_adaptor_2x2_0_output_01_waitrequest;        // adaptor_2x2_0:waiteRequest_01 -> mm_interconnect_1:adaptor_2x2_0_Output_01_waitrequest
	wire         mm_interconnect_1_adaptor_2x2_0_output_01_write;              // mm_interconnect_1:adaptor_2x2_0_Output_01_write -> adaptor_2x2_0:write_01
	wire   [7:0] mm_interconnect_1_adaptor_2x2_0_output_01_writedata;          // mm_interconnect_1:adaptor_2x2_0_Output_01_writedata -> adaptor_2x2_0:writeData_01
	wire         mm_interconnect_1_jtag_uart_01_avalon_jtag_slave_chipselect;  // mm_interconnect_1:jtag_uart_01_avalon_jtag_slave_chipselect -> jtag_uart_01:av_chipselect
	wire  [31:0] mm_interconnect_1_jtag_uart_01_avalon_jtag_slave_readdata;    // jtag_uart_01:av_readdata -> mm_interconnect_1:jtag_uart_01_avalon_jtag_slave_readdata
	wire         mm_interconnect_1_jtag_uart_01_avalon_jtag_slave_waitrequest; // jtag_uart_01:av_waitrequest -> mm_interconnect_1:jtag_uart_01_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_1_jtag_uart_01_avalon_jtag_slave_address;     // mm_interconnect_1:jtag_uart_01_avalon_jtag_slave_address -> jtag_uart_01:av_address
	wire         mm_interconnect_1_jtag_uart_01_avalon_jtag_slave_read;        // mm_interconnect_1:jtag_uart_01_avalon_jtag_slave_read -> jtag_uart_01:av_read_n
	wire         mm_interconnect_1_jtag_uart_01_avalon_jtag_slave_write;       // mm_interconnect_1:jtag_uart_01_avalon_jtag_slave_write -> jtag_uart_01:av_write_n
	wire  [31:0] mm_interconnect_1_jtag_uart_01_avalon_jtag_slave_writedata;   // mm_interconnect_1:jtag_uart_01_avalon_jtag_slave_writedata -> jtag_uart_01:av_writedata
	wire  [31:0] mm_interconnect_1_nios2_gen2_01_debug_mem_slave_readdata;     // nios2_gen2_01:debug_mem_slave_readdata -> mm_interconnect_1:nios2_gen2_01_debug_mem_slave_readdata
	wire         mm_interconnect_1_nios2_gen2_01_debug_mem_slave_waitrequest;  // nios2_gen2_01:debug_mem_slave_waitrequest -> mm_interconnect_1:nios2_gen2_01_debug_mem_slave_waitrequest
	wire         mm_interconnect_1_nios2_gen2_01_debug_mem_slave_debugaccess;  // mm_interconnect_1:nios2_gen2_01_debug_mem_slave_debugaccess -> nios2_gen2_01:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_1_nios2_gen2_01_debug_mem_slave_address;      // mm_interconnect_1:nios2_gen2_01_debug_mem_slave_address -> nios2_gen2_01:debug_mem_slave_address
	wire         mm_interconnect_1_nios2_gen2_01_debug_mem_slave_read;         // mm_interconnect_1:nios2_gen2_01_debug_mem_slave_read -> nios2_gen2_01:debug_mem_slave_read
	wire   [3:0] mm_interconnect_1_nios2_gen2_01_debug_mem_slave_byteenable;   // mm_interconnect_1:nios2_gen2_01_debug_mem_slave_byteenable -> nios2_gen2_01:debug_mem_slave_byteenable
	wire         mm_interconnect_1_nios2_gen2_01_debug_mem_slave_write;        // mm_interconnect_1:nios2_gen2_01_debug_mem_slave_write -> nios2_gen2_01:debug_mem_slave_write
	wire  [31:0] mm_interconnect_1_nios2_gen2_01_debug_mem_slave_writedata;    // mm_interconnect_1:nios2_gen2_01_debug_mem_slave_writedata -> nios2_gen2_01:debug_mem_slave_writedata
	wire         mm_interconnect_1_data_memory_01_s1_chipselect;               // mm_interconnect_1:Data_Memory_01_s1_chipselect -> Data_Memory_01:chipselect
	wire  [31:0] mm_interconnect_1_data_memory_01_s1_readdata;                 // Data_Memory_01:readdata -> mm_interconnect_1:Data_Memory_01_s1_readdata
	wire   [9:0] mm_interconnect_1_data_memory_01_s1_address;                  // mm_interconnect_1:Data_Memory_01_s1_address -> Data_Memory_01:address
	wire   [3:0] mm_interconnect_1_data_memory_01_s1_byteenable;               // mm_interconnect_1:Data_Memory_01_s1_byteenable -> Data_Memory_01:byteenable
	wire         mm_interconnect_1_data_memory_01_s1_write;                    // mm_interconnect_1:Data_Memory_01_s1_write -> Data_Memory_01:write
	wire  [31:0] mm_interconnect_1_data_memory_01_s1_writedata;                // mm_interconnect_1:Data_Memory_01_s1_writedata -> Data_Memory_01:writedata
	wire         mm_interconnect_1_data_memory_01_s1_clken;                    // mm_interconnect_1:Data_Memory_01_s1_clken -> Data_Memory_01:clken
	wire         mm_interconnect_1_instruction_memory_01_s1_chipselect;        // mm_interconnect_1:Instruction_Memory_01_s1_chipselect -> Instruction_Memory_01:chipselect
	wire  [31:0] mm_interconnect_1_instruction_memory_01_s1_readdata;          // Instruction_Memory_01:readdata -> mm_interconnect_1:Instruction_Memory_01_s1_readdata
	wire   [9:0] mm_interconnect_1_instruction_memory_01_s1_address;           // mm_interconnect_1:Instruction_Memory_01_s1_address -> Instruction_Memory_01:address
	wire   [3:0] mm_interconnect_1_instruction_memory_01_s1_byteenable;        // mm_interconnect_1:Instruction_Memory_01_s1_byteenable -> Instruction_Memory_01:byteenable
	wire         mm_interconnect_1_instruction_memory_01_s1_write;             // mm_interconnect_1:Instruction_Memory_01_s1_write -> Instruction_Memory_01:write
	wire  [31:0] mm_interconnect_1_instruction_memory_01_s1_writedata;         // mm_interconnect_1:Instruction_Memory_01_s1_writedata -> Instruction_Memory_01:writedata
	wire         mm_interconnect_1_instruction_memory_01_s1_clken;             // mm_interconnect_1:Instruction_Memory_01_s1_clken -> Instruction_Memory_01:clken
	wire  [31:0] nios2_gen2_10_data_master_readdata;                           // mm_interconnect_2:nios2_gen2_10_data_master_readdata -> nios2_gen2_10:d_readdata
	wire         nios2_gen2_10_data_master_waitrequest;                        // mm_interconnect_2:nios2_gen2_10_data_master_waitrequest -> nios2_gen2_10:d_waitrequest
	wire         nios2_gen2_10_data_master_debugaccess;                        // nios2_gen2_10:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_2:nios2_gen2_10_data_master_debugaccess
	wire  [13:0] nios2_gen2_10_data_master_address;                            // nios2_gen2_10:d_address -> mm_interconnect_2:nios2_gen2_10_data_master_address
	wire   [3:0] nios2_gen2_10_data_master_byteenable;                         // nios2_gen2_10:d_byteenable -> mm_interconnect_2:nios2_gen2_10_data_master_byteenable
	wire         nios2_gen2_10_data_master_read;                               // nios2_gen2_10:d_read -> mm_interconnect_2:nios2_gen2_10_data_master_read
	wire         nios2_gen2_10_data_master_write;                              // nios2_gen2_10:d_write -> mm_interconnect_2:nios2_gen2_10_data_master_write
	wire  [31:0] nios2_gen2_10_data_master_writedata;                          // nios2_gen2_10:d_writedata -> mm_interconnect_2:nios2_gen2_10_data_master_writedata
	wire  [31:0] nios2_gen2_10_instruction_master_readdata;                    // mm_interconnect_2:nios2_gen2_10_instruction_master_readdata -> nios2_gen2_10:i_readdata
	wire         nios2_gen2_10_instruction_master_waitrequest;                 // mm_interconnect_2:nios2_gen2_10_instruction_master_waitrequest -> nios2_gen2_10:i_waitrequest
	wire  [13:0] nios2_gen2_10_instruction_master_address;                     // nios2_gen2_10:i_address -> mm_interconnect_2:nios2_gen2_10_instruction_master_address
	wire         nios2_gen2_10_instruction_master_read;                        // nios2_gen2_10:i_read -> mm_interconnect_2:nios2_gen2_10_instruction_master_read
	wire   [7:0] mm_interconnect_2_adaptor_2x2_0_input_10_readdata;            // adaptor_2x2_0:reaData_10 -> mm_interconnect_2:adaptor_2x2_0_Input_10_readdata
	wire         mm_interconnect_2_adaptor_2x2_0_input_10_read;                // mm_interconnect_2:adaptor_2x2_0_Input_10_read -> adaptor_2x2_0:read_10
	wire         mm_interconnect_2_adaptor_2x2_0_output_10_waitrequest;        // adaptor_2x2_0:waiteRequest_10 -> mm_interconnect_2:adaptor_2x2_0_Output_10_waitrequest
	wire         mm_interconnect_2_adaptor_2x2_0_output_10_write;              // mm_interconnect_2:adaptor_2x2_0_Output_10_write -> adaptor_2x2_0:write_10
	wire   [7:0] mm_interconnect_2_adaptor_2x2_0_output_10_writedata;          // mm_interconnect_2:adaptor_2x2_0_Output_10_writedata -> adaptor_2x2_0:writeData_10
	wire         mm_interconnect_2_jtag_uart_10_avalon_jtag_slave_chipselect;  // mm_interconnect_2:jtag_uart_10_avalon_jtag_slave_chipselect -> jtag_uart_10:av_chipselect
	wire  [31:0] mm_interconnect_2_jtag_uart_10_avalon_jtag_slave_readdata;    // jtag_uart_10:av_readdata -> mm_interconnect_2:jtag_uart_10_avalon_jtag_slave_readdata
	wire         mm_interconnect_2_jtag_uart_10_avalon_jtag_slave_waitrequest; // jtag_uart_10:av_waitrequest -> mm_interconnect_2:jtag_uart_10_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_2_jtag_uart_10_avalon_jtag_slave_address;     // mm_interconnect_2:jtag_uart_10_avalon_jtag_slave_address -> jtag_uart_10:av_address
	wire         mm_interconnect_2_jtag_uart_10_avalon_jtag_slave_read;        // mm_interconnect_2:jtag_uart_10_avalon_jtag_slave_read -> jtag_uart_10:av_read_n
	wire         mm_interconnect_2_jtag_uart_10_avalon_jtag_slave_write;       // mm_interconnect_2:jtag_uart_10_avalon_jtag_slave_write -> jtag_uart_10:av_write_n
	wire  [31:0] mm_interconnect_2_jtag_uart_10_avalon_jtag_slave_writedata;   // mm_interconnect_2:jtag_uart_10_avalon_jtag_slave_writedata -> jtag_uart_10:av_writedata
	wire  [31:0] mm_interconnect_2_nios2_gen2_10_debug_mem_slave_readdata;     // nios2_gen2_10:debug_mem_slave_readdata -> mm_interconnect_2:nios2_gen2_10_debug_mem_slave_readdata
	wire         mm_interconnect_2_nios2_gen2_10_debug_mem_slave_waitrequest;  // nios2_gen2_10:debug_mem_slave_waitrequest -> mm_interconnect_2:nios2_gen2_10_debug_mem_slave_waitrequest
	wire         mm_interconnect_2_nios2_gen2_10_debug_mem_slave_debugaccess;  // mm_interconnect_2:nios2_gen2_10_debug_mem_slave_debugaccess -> nios2_gen2_10:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_2_nios2_gen2_10_debug_mem_slave_address;      // mm_interconnect_2:nios2_gen2_10_debug_mem_slave_address -> nios2_gen2_10:debug_mem_slave_address
	wire         mm_interconnect_2_nios2_gen2_10_debug_mem_slave_read;         // mm_interconnect_2:nios2_gen2_10_debug_mem_slave_read -> nios2_gen2_10:debug_mem_slave_read
	wire   [3:0] mm_interconnect_2_nios2_gen2_10_debug_mem_slave_byteenable;   // mm_interconnect_2:nios2_gen2_10_debug_mem_slave_byteenable -> nios2_gen2_10:debug_mem_slave_byteenable
	wire         mm_interconnect_2_nios2_gen2_10_debug_mem_slave_write;        // mm_interconnect_2:nios2_gen2_10_debug_mem_slave_write -> nios2_gen2_10:debug_mem_slave_write
	wire  [31:0] mm_interconnect_2_nios2_gen2_10_debug_mem_slave_writedata;    // mm_interconnect_2:nios2_gen2_10_debug_mem_slave_writedata -> nios2_gen2_10:debug_mem_slave_writedata
	wire         mm_interconnect_2_data_memory_10_s1_chipselect;               // mm_interconnect_2:Data_Memory_10_s1_chipselect -> Data_Memory_10:chipselect
	wire  [31:0] mm_interconnect_2_data_memory_10_s1_readdata;                 // Data_Memory_10:readdata -> mm_interconnect_2:Data_Memory_10_s1_readdata
	wire   [9:0] mm_interconnect_2_data_memory_10_s1_address;                  // mm_interconnect_2:Data_Memory_10_s1_address -> Data_Memory_10:address
	wire   [3:0] mm_interconnect_2_data_memory_10_s1_byteenable;               // mm_interconnect_2:Data_Memory_10_s1_byteenable -> Data_Memory_10:byteenable
	wire         mm_interconnect_2_data_memory_10_s1_write;                    // mm_interconnect_2:Data_Memory_10_s1_write -> Data_Memory_10:write
	wire  [31:0] mm_interconnect_2_data_memory_10_s1_writedata;                // mm_interconnect_2:Data_Memory_10_s1_writedata -> Data_Memory_10:writedata
	wire         mm_interconnect_2_data_memory_10_s1_clken;                    // mm_interconnect_2:Data_Memory_10_s1_clken -> Data_Memory_10:clken
	wire         mm_interconnect_2_instruction_memory_10_s1_chipselect;        // mm_interconnect_2:Instruction_Memory_10_s1_chipselect -> Instruction_Memory_10:chipselect
	wire  [31:0] mm_interconnect_2_instruction_memory_10_s1_readdata;          // Instruction_Memory_10:readdata -> mm_interconnect_2:Instruction_Memory_10_s1_readdata
	wire   [9:0] mm_interconnect_2_instruction_memory_10_s1_address;           // mm_interconnect_2:Instruction_Memory_10_s1_address -> Instruction_Memory_10:address
	wire   [3:0] mm_interconnect_2_instruction_memory_10_s1_byteenable;        // mm_interconnect_2:Instruction_Memory_10_s1_byteenable -> Instruction_Memory_10:byteenable
	wire         mm_interconnect_2_instruction_memory_10_s1_write;             // mm_interconnect_2:Instruction_Memory_10_s1_write -> Instruction_Memory_10:write
	wire  [31:0] mm_interconnect_2_instruction_memory_10_s1_writedata;         // mm_interconnect_2:Instruction_Memory_10_s1_writedata -> Instruction_Memory_10:writedata
	wire         mm_interconnect_2_instruction_memory_10_s1_clken;             // mm_interconnect_2:Instruction_Memory_10_s1_clken -> Instruction_Memory_10:clken
	wire  [31:0] nios2_gen2_11_data_master_readdata;                           // mm_interconnect_3:nios2_gen2_11_data_master_readdata -> nios2_gen2_11:d_readdata
	wire         nios2_gen2_11_data_master_waitrequest;                        // mm_interconnect_3:nios2_gen2_11_data_master_waitrequest -> nios2_gen2_11:d_waitrequest
	wire         nios2_gen2_11_data_master_debugaccess;                        // nios2_gen2_11:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_3:nios2_gen2_11_data_master_debugaccess
	wire  [13:0] nios2_gen2_11_data_master_address;                            // nios2_gen2_11:d_address -> mm_interconnect_3:nios2_gen2_11_data_master_address
	wire   [3:0] nios2_gen2_11_data_master_byteenable;                         // nios2_gen2_11:d_byteenable -> mm_interconnect_3:nios2_gen2_11_data_master_byteenable
	wire         nios2_gen2_11_data_master_read;                               // nios2_gen2_11:d_read -> mm_interconnect_3:nios2_gen2_11_data_master_read
	wire         nios2_gen2_11_data_master_write;                              // nios2_gen2_11:d_write -> mm_interconnect_3:nios2_gen2_11_data_master_write
	wire  [31:0] nios2_gen2_11_data_master_writedata;                          // nios2_gen2_11:d_writedata -> mm_interconnect_3:nios2_gen2_11_data_master_writedata
	wire  [31:0] nios2_gen2_11_instruction_master_readdata;                    // mm_interconnect_3:nios2_gen2_11_instruction_master_readdata -> nios2_gen2_11:i_readdata
	wire         nios2_gen2_11_instruction_master_waitrequest;                 // mm_interconnect_3:nios2_gen2_11_instruction_master_waitrequest -> nios2_gen2_11:i_waitrequest
	wire  [13:0] nios2_gen2_11_instruction_master_address;                     // nios2_gen2_11:i_address -> mm_interconnect_3:nios2_gen2_11_instruction_master_address
	wire         nios2_gen2_11_instruction_master_read;                        // nios2_gen2_11:i_read -> mm_interconnect_3:nios2_gen2_11_instruction_master_read
	wire   [7:0] mm_interconnect_3_adaptor_2x2_0_input_11_readdata;            // adaptor_2x2_0:reaData_11 -> mm_interconnect_3:adaptor_2x2_0_Input_11_readdata
	wire         mm_interconnect_3_adaptor_2x2_0_input_11_read;                // mm_interconnect_3:adaptor_2x2_0_Input_11_read -> adaptor_2x2_0:read_11
	wire         mm_interconnect_3_adaptor_2x2_0_output_11_waitrequest;        // adaptor_2x2_0:waiteRequest_11 -> mm_interconnect_3:adaptor_2x2_0_Output_11_waitrequest
	wire         mm_interconnect_3_adaptor_2x2_0_output_11_write;              // mm_interconnect_3:adaptor_2x2_0_Output_11_write -> adaptor_2x2_0:write_11
	wire   [7:0] mm_interconnect_3_adaptor_2x2_0_output_11_writedata;          // mm_interconnect_3:adaptor_2x2_0_Output_11_writedata -> adaptor_2x2_0:writeData_11
	wire         mm_interconnect_3_jtag_uart_11_avalon_jtag_slave_chipselect;  // mm_interconnect_3:jtag_uart_11_avalon_jtag_slave_chipselect -> jtag_uart_11:av_chipselect
	wire  [31:0] mm_interconnect_3_jtag_uart_11_avalon_jtag_slave_readdata;    // jtag_uart_11:av_readdata -> mm_interconnect_3:jtag_uart_11_avalon_jtag_slave_readdata
	wire         mm_interconnect_3_jtag_uart_11_avalon_jtag_slave_waitrequest; // jtag_uart_11:av_waitrequest -> mm_interconnect_3:jtag_uart_11_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_3_jtag_uart_11_avalon_jtag_slave_address;     // mm_interconnect_3:jtag_uart_11_avalon_jtag_slave_address -> jtag_uart_11:av_address
	wire         mm_interconnect_3_jtag_uart_11_avalon_jtag_slave_read;        // mm_interconnect_3:jtag_uart_11_avalon_jtag_slave_read -> jtag_uart_11:av_read_n
	wire         mm_interconnect_3_jtag_uart_11_avalon_jtag_slave_write;       // mm_interconnect_3:jtag_uart_11_avalon_jtag_slave_write -> jtag_uart_11:av_write_n
	wire  [31:0] mm_interconnect_3_jtag_uart_11_avalon_jtag_slave_writedata;   // mm_interconnect_3:jtag_uart_11_avalon_jtag_slave_writedata -> jtag_uart_11:av_writedata
	wire  [31:0] mm_interconnect_3_nios2_gen2_11_debug_mem_slave_readdata;     // nios2_gen2_11:debug_mem_slave_readdata -> mm_interconnect_3:nios2_gen2_11_debug_mem_slave_readdata
	wire         mm_interconnect_3_nios2_gen2_11_debug_mem_slave_waitrequest;  // nios2_gen2_11:debug_mem_slave_waitrequest -> mm_interconnect_3:nios2_gen2_11_debug_mem_slave_waitrequest
	wire         mm_interconnect_3_nios2_gen2_11_debug_mem_slave_debugaccess;  // mm_interconnect_3:nios2_gen2_11_debug_mem_slave_debugaccess -> nios2_gen2_11:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_3_nios2_gen2_11_debug_mem_slave_address;      // mm_interconnect_3:nios2_gen2_11_debug_mem_slave_address -> nios2_gen2_11:debug_mem_slave_address
	wire         mm_interconnect_3_nios2_gen2_11_debug_mem_slave_read;         // mm_interconnect_3:nios2_gen2_11_debug_mem_slave_read -> nios2_gen2_11:debug_mem_slave_read
	wire   [3:0] mm_interconnect_3_nios2_gen2_11_debug_mem_slave_byteenable;   // mm_interconnect_3:nios2_gen2_11_debug_mem_slave_byteenable -> nios2_gen2_11:debug_mem_slave_byteenable
	wire         mm_interconnect_3_nios2_gen2_11_debug_mem_slave_write;        // mm_interconnect_3:nios2_gen2_11_debug_mem_slave_write -> nios2_gen2_11:debug_mem_slave_write
	wire  [31:0] mm_interconnect_3_nios2_gen2_11_debug_mem_slave_writedata;    // mm_interconnect_3:nios2_gen2_11_debug_mem_slave_writedata -> nios2_gen2_11:debug_mem_slave_writedata
	wire         mm_interconnect_3_data_memory_11_s1_chipselect;               // mm_interconnect_3:Data_Memory_11_s1_chipselect -> Data_Memory_11:chipselect
	wire  [31:0] mm_interconnect_3_data_memory_11_s1_readdata;                 // Data_Memory_11:readdata -> mm_interconnect_3:Data_Memory_11_s1_readdata
	wire   [9:0] mm_interconnect_3_data_memory_11_s1_address;                  // mm_interconnect_3:Data_Memory_11_s1_address -> Data_Memory_11:address
	wire   [3:0] mm_interconnect_3_data_memory_11_s1_byteenable;               // mm_interconnect_3:Data_Memory_11_s1_byteenable -> Data_Memory_11:byteenable
	wire         mm_interconnect_3_data_memory_11_s1_write;                    // mm_interconnect_3:Data_Memory_11_s1_write -> Data_Memory_11:write
	wire  [31:0] mm_interconnect_3_data_memory_11_s1_writedata;                // mm_interconnect_3:Data_Memory_11_s1_writedata -> Data_Memory_11:writedata
	wire         mm_interconnect_3_data_memory_11_s1_clken;                    // mm_interconnect_3:Data_Memory_11_s1_clken -> Data_Memory_11:clken
	wire         mm_interconnect_3_instruction_memory_11_s1_chipselect;        // mm_interconnect_3:Instruction_Memory_11_s1_chipselect -> Instruction_Memory_11:chipselect
	wire  [31:0] mm_interconnect_3_instruction_memory_11_s1_readdata;          // Instruction_Memory_11:readdata -> mm_interconnect_3:Instruction_Memory_11_s1_readdata
	wire   [9:0] mm_interconnect_3_instruction_memory_11_s1_address;           // mm_interconnect_3:Instruction_Memory_11_s1_address -> Instruction_Memory_11:address
	wire   [3:0] mm_interconnect_3_instruction_memory_11_s1_byteenable;        // mm_interconnect_3:Instruction_Memory_11_s1_byteenable -> Instruction_Memory_11:byteenable
	wire         mm_interconnect_3_instruction_memory_11_s1_write;             // mm_interconnect_3:Instruction_Memory_11_s1_write -> Instruction_Memory_11:write
	wire  [31:0] mm_interconnect_3_instruction_memory_11_s1_writedata;         // mm_interconnect_3:Instruction_Memory_11_s1_writedata -> Instruction_Memory_11:writedata
	wire         mm_interconnect_3_instruction_memory_11_s1_clken;             // mm_interconnect_3:Instruction_Memory_11_s1_clken -> Instruction_Memory_11:clken
	wire         irq_mapper_receiver0_irq;                                     // adaptor_2x2_0:irq_00 -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                     // jtag_uart_00:av_irq -> irq_mapper:receiver1_irq
	wire  [31:0] nios2_gen2_00_irq_irq;                                        // irq_mapper:sender_irq -> nios2_gen2_00:irq
	wire         irq_mapper_001_receiver0_irq;                                 // adaptor_2x2_0:irq_01 -> irq_mapper_001:receiver0_irq
	wire         irq_mapper_001_receiver1_irq;                                 // jtag_uart_01:av_irq -> irq_mapper_001:receiver1_irq
	wire  [31:0] nios2_gen2_01_irq_irq;                                        // irq_mapper_001:sender_irq -> nios2_gen2_01:irq
	wire         irq_mapper_002_receiver0_irq;                                 // adaptor_2x2_0:irq_10 -> irq_mapper_002:receiver0_irq
	wire         irq_mapper_002_receiver1_irq;                                 // jtag_uart_10:av_irq -> irq_mapper_002:receiver1_irq
	wire  [31:0] nios2_gen2_10_irq_irq;                                        // irq_mapper_002:sender_irq -> nios2_gen2_10:irq
	wire         irq_mapper_003_receiver0_irq;                                 // adaptor_2x2_0:irq_11 -> irq_mapper_003:receiver0_irq
	wire         irq_mapper_003_receiver1_irq;                                 // jtag_uart_11:av_irq -> irq_mapper_003:receiver1_irq
	wire  [31:0] nios2_gen2_11_irq_irq;                                        // irq_mapper_003:sender_irq -> nios2_gen2_11:irq
	wire         rst_controller_reset_out_reset;                               // rst_controller:reset_out -> [Data_Memory_00:reset, Data_Memory_01:reset, Data_Memory_10:reset, Data_Memory_11:reset, Instruction_Memory_00:reset, Instruction_Memory_01:reset, Instruction_Memory_10:reset, Instruction_Memory_11:reset, adaptor_2x2_0:reset, irq_mapper:reset, irq_mapper_001:reset, irq_mapper_002:reset, irq_mapper_003:reset, jtag_uart_00:rst_n, jtag_uart_01:rst_n, jtag_uart_10:rst_n, jtag_uart_11:rst_n, mm_interconnect_0:nios2_gen2_00_reset_reset_bridge_in_reset_reset, mm_interconnect_1:nios2_gen2_01_reset_reset_bridge_in_reset_reset, mm_interconnect_2:nios2_gen2_10_reset_reset_bridge_in_reset_reset, mm_interconnect_3:nios2_gen2_11_reset_reset_bridge_in_reset_reset, nios2_gen2_00:reset_n, nios2_gen2_01:reset_n, nios2_gen2_10:reset_n, nios2_gen2_11:reset_n, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                           // rst_controller:reset_req -> [Data_Memory_00:reset_req, Data_Memory_01:reset_req, Data_Memory_10:reset_req, Data_Memory_11:reset_req, Instruction_Memory_00:reset_req, Instruction_Memory_01:reset_req, Instruction_Memory_10:reset_req, Instruction_Memory_11:reset_req, nios2_gen2_00:reset_req, nios2_gen2_01:reset_req, nios2_gen2_10:reset_req, nios2_gen2_11:reset_req, rst_translator:reset_req_in]

	adaptor2x2_Data_Memory_00 data_memory_00 (
		.clk        (clk_clk),                                        //   clk1.clk
		.address    (mm_interconnect_0_data_memory_00_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_data_memory_00_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_data_memory_00_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_data_memory_00_s1_write),      //       .write
		.readdata   (mm_interconnect_0_data_memory_00_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_data_memory_00_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_data_memory_00_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                 // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),             //       .reset_req
		.freeze     (1'b0)                                            // (terminated)
	);

	adaptor2x2_Data_Memory_01 data_memory_01 (
		.clk        (clk_clk),                                        //   clk1.clk
		.address    (mm_interconnect_1_data_memory_01_s1_address),    //     s1.address
		.clken      (mm_interconnect_1_data_memory_01_s1_clken),      //       .clken
		.chipselect (mm_interconnect_1_data_memory_01_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_1_data_memory_01_s1_write),      //       .write
		.readdata   (mm_interconnect_1_data_memory_01_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_1_data_memory_01_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_1_data_memory_01_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                 // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),             //       .reset_req
		.freeze     (1'b0)                                            // (terminated)
	);

	adaptor2x2_Data_Memory_10 data_memory_10 (
		.clk        (clk_clk),                                        //   clk1.clk
		.address    (mm_interconnect_2_data_memory_10_s1_address),    //     s1.address
		.clken      (mm_interconnect_2_data_memory_10_s1_clken),      //       .clken
		.chipselect (mm_interconnect_2_data_memory_10_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_2_data_memory_10_s1_write),      //       .write
		.readdata   (mm_interconnect_2_data_memory_10_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_2_data_memory_10_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_2_data_memory_10_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                 // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),             //       .reset_req
		.freeze     (1'b0)                                            // (terminated)
	);

	adaptor2x2_Data_Memory_11 data_memory_11 (
		.clk        (clk_clk),                                        //   clk1.clk
		.address    (mm_interconnect_3_data_memory_11_s1_address),    //     s1.address
		.clken      (mm_interconnect_3_data_memory_11_s1_clken),      //       .clken
		.chipselect (mm_interconnect_3_data_memory_11_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_3_data_memory_11_s1_write),      //       .write
		.readdata   (mm_interconnect_3_data_memory_11_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_3_data_memory_11_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_3_data_memory_11_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                 // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),             //       .reset_req
		.freeze     (1'b0)                                            // (terminated)
	);

	adaptor2x2_Instruction_Memory_00 instruction_memory_00 (
		.clk        (clk_clk),                                               //   clk1.clk
		.address    (mm_interconnect_0_instruction_memory_00_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_instruction_memory_00_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_instruction_memory_00_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_instruction_memory_00_s1_write),      //       .write
		.readdata   (mm_interconnect_0_instruction_memory_00_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_instruction_memory_00_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_instruction_memory_00_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                        // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),                    //       .reset_req
		.freeze     (1'b0)                                                   // (terminated)
	);

	adaptor2x2_Instruction_Memory_01 instruction_memory_01 (
		.clk        (clk_clk),                                               //   clk1.clk
		.address    (mm_interconnect_1_instruction_memory_01_s1_address),    //     s1.address
		.clken      (mm_interconnect_1_instruction_memory_01_s1_clken),      //       .clken
		.chipselect (mm_interconnect_1_instruction_memory_01_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_1_instruction_memory_01_s1_write),      //       .write
		.readdata   (mm_interconnect_1_instruction_memory_01_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_1_instruction_memory_01_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_1_instruction_memory_01_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                        // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),                    //       .reset_req
		.freeze     (1'b0)                                                   // (terminated)
	);

	adaptor2x2_Instruction_Memory_10 instruction_memory_10 (
		.clk        (clk_clk),                                               //   clk1.clk
		.address    (mm_interconnect_2_instruction_memory_10_s1_address),    //     s1.address
		.clken      (mm_interconnect_2_instruction_memory_10_s1_clken),      //       .clken
		.chipselect (mm_interconnect_2_instruction_memory_10_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_2_instruction_memory_10_s1_write),      //       .write
		.readdata   (mm_interconnect_2_instruction_memory_10_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_2_instruction_memory_10_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_2_instruction_memory_10_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                        // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),                    //       .reset_req
		.freeze     (1'b0)                                                   // (terminated)
	);

	adaptor2x2_Instruction_Memory_11 instruction_memory_11 (
		.clk        (clk_clk),                                               //   clk1.clk
		.address    (mm_interconnect_3_instruction_memory_11_s1_address),    //     s1.address
		.clken      (mm_interconnect_3_instruction_memory_11_s1_clken),      //       .clken
		.chipselect (mm_interconnect_3_instruction_memory_11_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_3_instruction_memory_11_s1_write),      //       .write
		.readdata   (mm_interconnect_3_instruction_memory_11_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_3_instruction_memory_11_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_3_instruction_memory_11_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                        // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),                    //       .reset_req
		.freeze     (1'b0)                                                   // (terminated)
	);

	adaptor #(
		.DataWidth (8)
	) adaptor_2x2_0 (
		.clock           (clk_clk),                                               //          clock_sink.clk
		.reset           (rst_controller_reset_out_reset),                        //          reset_sink.reset
		.reaData_00      (mm_interconnect_0_adaptor_2x2_0_input_00_readdata),     //            Input_00.readdata
		.read_00         (mm_interconnect_0_adaptor_2x2_0_input_00_read),         //                    .read
		.reaData_01      (mm_interconnect_1_adaptor_2x2_0_input_01_readdata),     //            Input_01.readdata
		.read_01         (mm_interconnect_1_adaptor_2x2_0_input_01_read),         //                    .read
		.read_10         (mm_interconnect_2_adaptor_2x2_0_input_10_read),         //            Input_10.read
		.reaData_10      (mm_interconnect_2_adaptor_2x2_0_input_10_readdata),     //                    .readdata
		.reaData_11      (mm_interconnect_3_adaptor_2x2_0_input_11_readdata),     //            Input_11.readdata
		.read_11         (mm_interconnect_3_adaptor_2x2_0_input_11_read),         //                    .read
		.writeData_00    (mm_interconnect_0_adaptor_2x2_0_output_00_writedata),   //           Output_00.writedata
		.write_00        (mm_interconnect_0_adaptor_2x2_0_output_00_write),       //                    .write
		.waiteRequest_00 (mm_interconnect_0_adaptor_2x2_0_output_00_waitrequest), //                    .waitrequest
		.writeData_01    (mm_interconnect_1_adaptor_2x2_0_output_01_writedata),   //           Output_01.writedata
		.write_01        (mm_interconnect_1_adaptor_2x2_0_output_01_write),       //                    .write
		.waiteRequest_01 (mm_interconnect_1_adaptor_2x2_0_output_01_waitrequest), //                    .waitrequest
		.writeData_10    (mm_interconnect_2_adaptor_2x2_0_output_10_writedata),   //           Output_10.writedata
		.write_10        (mm_interconnect_2_adaptor_2x2_0_output_10_write),       //                    .write
		.waiteRequest_10 (mm_interconnect_2_adaptor_2x2_0_output_10_waitrequest), //                    .waitrequest
		.writeData_11    (mm_interconnect_3_adaptor_2x2_0_output_11_writedata),   //           Output_11.writedata
		.write_11        (mm_interconnect_3_adaptor_2x2_0_output_11_write),       //                    .write
		.waiteRequest_11 (mm_interconnect_3_adaptor_2x2_0_output_11_waitrequest), //                    .waitrequest
		.irq_00          (irq_mapper_receiver0_irq),                              // interrupt_sender_00.irq
		.irq_01          (irq_mapper_001_receiver0_irq),                          // interrupt_sender_01.irq
		.irq_10          (irq_mapper_002_receiver0_irq),                          // interrupt_sender_10.irq
		.irq_11          (irq_mapper_003_receiver0_irq)                           // interrupt_sender_11.irq
	);

	adaptor2x2_jtag_uart_00 jtag_uart_00 (
		.clk            (clk_clk),                                                      //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                              //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_00_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_00_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_00_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_00_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_00_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_00_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_00_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                      //               irq.irq
	);

	adaptor2x2_jtag_uart_00 jtag_uart_01 (
		.clk            (clk_clk),                                                      //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                              //             reset.reset_n
		.av_chipselect  (mm_interconnect_1_jtag_uart_01_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_1_jtag_uart_01_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_1_jtag_uart_01_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_1_jtag_uart_01_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_1_jtag_uart_01_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_1_jtag_uart_01_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_1_jtag_uart_01_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_001_receiver1_irq)                                  //               irq.irq
	);

	adaptor2x2_jtag_uart_00 jtag_uart_10 (
		.clk            (clk_clk),                                                      //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                              //             reset.reset_n
		.av_chipselect  (mm_interconnect_2_jtag_uart_10_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_2_jtag_uart_10_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_2_jtag_uart_10_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_2_jtag_uart_10_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_2_jtag_uart_10_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_2_jtag_uart_10_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_2_jtag_uart_10_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_002_receiver1_irq)                                  //               irq.irq
	);

	adaptor2x2_jtag_uart_00 jtag_uart_11 (
		.clk            (clk_clk),                                                      //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                              //             reset.reset_n
		.av_chipselect  (mm_interconnect_3_jtag_uart_11_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_3_jtag_uart_11_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_3_jtag_uart_11_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_3_jtag_uart_11_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_3_jtag_uart_11_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_3_jtag_uart_11_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_3_jtag_uart_11_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_003_receiver1_irq)                                  //               irq.irq
	);

	adaptor2x2_nios2_gen2_00 nios2_gen2_00 (
		.clk                                 (clk_clk),                                                     //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                             //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                          //                          .reset_req
		.d_address                           (nios2_gen2_00_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_00_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_00_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_00_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_00_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_00_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_00_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_00_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_00_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_00_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_00_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_00_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_gen2_00_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                            //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_00_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_00_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_00_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_00_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_00_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_00_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_00_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_00_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                             // custom_instruction_master.readra
	);

	adaptor2x2_nios2_gen2_01 nios2_gen2_01 (
		.clk                                 (clk_clk),                                                     //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                             //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                          //                          .reset_req
		.d_address                           (nios2_gen2_01_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_01_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_01_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_01_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_01_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_01_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_01_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_01_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_01_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_01_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_01_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_01_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_gen2_01_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                            //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_1_nios2_gen2_01_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_1_nios2_gen2_01_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_1_nios2_gen2_01_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_1_nios2_gen2_01_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_1_nios2_gen2_01_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_1_nios2_gen2_01_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_1_nios2_gen2_01_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_1_nios2_gen2_01_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                             // custom_instruction_master.readra
	);

	adaptor2x2_nios2_gen2_10 nios2_gen2_10 (
		.clk                                 (clk_clk),                                                     //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                             //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                          //                          .reset_req
		.d_address                           (nios2_gen2_10_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_10_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_10_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_10_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_10_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_10_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_10_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_10_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_10_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_10_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_10_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_10_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_gen2_10_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                            //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_2_nios2_gen2_10_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_2_nios2_gen2_10_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_2_nios2_gen2_10_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_2_nios2_gen2_10_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_2_nios2_gen2_10_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_2_nios2_gen2_10_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_2_nios2_gen2_10_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_2_nios2_gen2_10_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                             // custom_instruction_master.readra
	);

	adaptor2x2_nios2_gen2_11 nios2_gen2_11 (
		.clk                                 (clk_clk),                                                     //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                             //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                          //                          .reset_req
		.d_address                           (nios2_gen2_11_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_11_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_11_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_11_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_11_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_11_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_11_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_11_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_11_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_11_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_11_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_11_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_gen2_11_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                            //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_3_nios2_gen2_11_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_3_nios2_gen2_11_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_3_nios2_gen2_11_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_3_nios2_gen2_11_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_3_nios2_gen2_11_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_3_nios2_gen2_11_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_3_nios2_gen2_11_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_3_nios2_gen2_11_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                             // custom_instruction_master.readra
	);

	adaptor2x2_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                   (clk_clk),                                                      //                                 clk_0_clk.clk
		.nios2_gen2_00_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                               // nios2_gen2_00_reset_reset_bridge_in_reset.reset
		.nios2_gen2_00_data_master_address               (nios2_gen2_00_data_master_address),                            //                 nios2_gen2_00_data_master.address
		.nios2_gen2_00_data_master_waitrequest           (nios2_gen2_00_data_master_waitrequest),                        //                                          .waitrequest
		.nios2_gen2_00_data_master_byteenable            (nios2_gen2_00_data_master_byteenable),                         //                                          .byteenable
		.nios2_gen2_00_data_master_read                  (nios2_gen2_00_data_master_read),                               //                                          .read
		.nios2_gen2_00_data_master_readdata              (nios2_gen2_00_data_master_readdata),                           //                                          .readdata
		.nios2_gen2_00_data_master_write                 (nios2_gen2_00_data_master_write),                              //                                          .write
		.nios2_gen2_00_data_master_writedata             (nios2_gen2_00_data_master_writedata),                          //                                          .writedata
		.nios2_gen2_00_data_master_debugaccess           (nios2_gen2_00_data_master_debugaccess),                        //                                          .debugaccess
		.nios2_gen2_00_instruction_master_address        (nios2_gen2_00_instruction_master_address),                     //          nios2_gen2_00_instruction_master.address
		.nios2_gen2_00_instruction_master_waitrequest    (nios2_gen2_00_instruction_master_waitrequest),                 //                                          .waitrequest
		.nios2_gen2_00_instruction_master_read           (nios2_gen2_00_instruction_master_read),                        //                                          .read
		.nios2_gen2_00_instruction_master_readdata       (nios2_gen2_00_instruction_master_readdata),                    //                                          .readdata
		.adaptor_2x2_0_Input_00_read                     (mm_interconnect_0_adaptor_2x2_0_input_00_read),                //                    adaptor_2x2_0_Input_00.read
		.adaptor_2x2_0_Input_00_readdata                 (mm_interconnect_0_adaptor_2x2_0_input_00_readdata),            //                                          .readdata
		.adaptor_2x2_0_Output_00_write                   (mm_interconnect_0_adaptor_2x2_0_output_00_write),              //                   adaptor_2x2_0_Output_00.write
		.adaptor_2x2_0_Output_00_writedata               (mm_interconnect_0_adaptor_2x2_0_output_00_writedata),          //                                          .writedata
		.adaptor_2x2_0_Output_00_waitrequest             (mm_interconnect_0_adaptor_2x2_0_output_00_waitrequest),        //                                          .waitrequest
		.Data_Memory_00_s1_address                       (mm_interconnect_0_data_memory_00_s1_address),                  //                         Data_Memory_00_s1.address
		.Data_Memory_00_s1_write                         (mm_interconnect_0_data_memory_00_s1_write),                    //                                          .write
		.Data_Memory_00_s1_readdata                      (mm_interconnect_0_data_memory_00_s1_readdata),                 //                                          .readdata
		.Data_Memory_00_s1_writedata                     (mm_interconnect_0_data_memory_00_s1_writedata),                //                                          .writedata
		.Data_Memory_00_s1_byteenable                    (mm_interconnect_0_data_memory_00_s1_byteenable),               //                                          .byteenable
		.Data_Memory_00_s1_chipselect                    (mm_interconnect_0_data_memory_00_s1_chipselect),               //                                          .chipselect
		.Data_Memory_00_s1_clken                         (mm_interconnect_0_data_memory_00_s1_clken),                    //                                          .clken
		.Instruction_Memory_00_s1_address                (mm_interconnect_0_instruction_memory_00_s1_address),           //                  Instruction_Memory_00_s1.address
		.Instruction_Memory_00_s1_write                  (mm_interconnect_0_instruction_memory_00_s1_write),             //                                          .write
		.Instruction_Memory_00_s1_readdata               (mm_interconnect_0_instruction_memory_00_s1_readdata),          //                                          .readdata
		.Instruction_Memory_00_s1_writedata              (mm_interconnect_0_instruction_memory_00_s1_writedata),         //                                          .writedata
		.Instruction_Memory_00_s1_byteenable             (mm_interconnect_0_instruction_memory_00_s1_byteenable),        //                                          .byteenable
		.Instruction_Memory_00_s1_chipselect             (mm_interconnect_0_instruction_memory_00_s1_chipselect),        //                                          .chipselect
		.Instruction_Memory_00_s1_clken                  (mm_interconnect_0_instruction_memory_00_s1_clken),             //                                          .clken
		.jtag_uart_00_avalon_jtag_slave_address          (mm_interconnect_0_jtag_uart_00_avalon_jtag_slave_address),     //            jtag_uart_00_avalon_jtag_slave.address
		.jtag_uart_00_avalon_jtag_slave_write            (mm_interconnect_0_jtag_uart_00_avalon_jtag_slave_write),       //                                          .write
		.jtag_uart_00_avalon_jtag_slave_read             (mm_interconnect_0_jtag_uart_00_avalon_jtag_slave_read),        //                                          .read
		.jtag_uart_00_avalon_jtag_slave_readdata         (mm_interconnect_0_jtag_uart_00_avalon_jtag_slave_readdata),    //                                          .readdata
		.jtag_uart_00_avalon_jtag_slave_writedata        (mm_interconnect_0_jtag_uart_00_avalon_jtag_slave_writedata),   //                                          .writedata
		.jtag_uart_00_avalon_jtag_slave_waitrequest      (mm_interconnect_0_jtag_uart_00_avalon_jtag_slave_waitrequest), //                                          .waitrequest
		.jtag_uart_00_avalon_jtag_slave_chipselect       (mm_interconnect_0_jtag_uart_00_avalon_jtag_slave_chipselect),  //                                          .chipselect
		.nios2_gen2_00_debug_mem_slave_address           (mm_interconnect_0_nios2_gen2_00_debug_mem_slave_address),      //             nios2_gen2_00_debug_mem_slave.address
		.nios2_gen2_00_debug_mem_slave_write             (mm_interconnect_0_nios2_gen2_00_debug_mem_slave_write),        //                                          .write
		.nios2_gen2_00_debug_mem_slave_read              (mm_interconnect_0_nios2_gen2_00_debug_mem_slave_read),         //                                          .read
		.nios2_gen2_00_debug_mem_slave_readdata          (mm_interconnect_0_nios2_gen2_00_debug_mem_slave_readdata),     //                                          .readdata
		.nios2_gen2_00_debug_mem_slave_writedata         (mm_interconnect_0_nios2_gen2_00_debug_mem_slave_writedata),    //                                          .writedata
		.nios2_gen2_00_debug_mem_slave_byteenable        (mm_interconnect_0_nios2_gen2_00_debug_mem_slave_byteenable),   //                                          .byteenable
		.nios2_gen2_00_debug_mem_slave_waitrequest       (mm_interconnect_0_nios2_gen2_00_debug_mem_slave_waitrequest),  //                                          .waitrequest
		.nios2_gen2_00_debug_mem_slave_debugaccess       (mm_interconnect_0_nios2_gen2_00_debug_mem_slave_debugaccess)   //                                          .debugaccess
	);

	adaptor2x2_mm_interconnect_1 mm_interconnect_1 (
		.clk_0_clk_clk                                   (clk_clk),                                                      //                                 clk_0_clk.clk
		.nios2_gen2_01_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                               // nios2_gen2_01_reset_reset_bridge_in_reset.reset
		.nios2_gen2_01_data_master_address               (nios2_gen2_01_data_master_address),                            //                 nios2_gen2_01_data_master.address
		.nios2_gen2_01_data_master_waitrequest           (nios2_gen2_01_data_master_waitrequest),                        //                                          .waitrequest
		.nios2_gen2_01_data_master_byteenable            (nios2_gen2_01_data_master_byteenable),                         //                                          .byteenable
		.nios2_gen2_01_data_master_read                  (nios2_gen2_01_data_master_read),                               //                                          .read
		.nios2_gen2_01_data_master_readdata              (nios2_gen2_01_data_master_readdata),                           //                                          .readdata
		.nios2_gen2_01_data_master_write                 (nios2_gen2_01_data_master_write),                              //                                          .write
		.nios2_gen2_01_data_master_writedata             (nios2_gen2_01_data_master_writedata),                          //                                          .writedata
		.nios2_gen2_01_data_master_debugaccess           (nios2_gen2_01_data_master_debugaccess),                        //                                          .debugaccess
		.nios2_gen2_01_instruction_master_address        (nios2_gen2_01_instruction_master_address),                     //          nios2_gen2_01_instruction_master.address
		.nios2_gen2_01_instruction_master_waitrequest    (nios2_gen2_01_instruction_master_waitrequest),                 //                                          .waitrequest
		.nios2_gen2_01_instruction_master_read           (nios2_gen2_01_instruction_master_read),                        //                                          .read
		.nios2_gen2_01_instruction_master_readdata       (nios2_gen2_01_instruction_master_readdata),                    //                                          .readdata
		.adaptor_2x2_0_Input_01_read                     (mm_interconnect_1_adaptor_2x2_0_input_01_read),                //                    adaptor_2x2_0_Input_01.read
		.adaptor_2x2_0_Input_01_readdata                 (mm_interconnect_1_adaptor_2x2_0_input_01_readdata),            //                                          .readdata
		.adaptor_2x2_0_Output_01_write                   (mm_interconnect_1_adaptor_2x2_0_output_01_write),              //                   adaptor_2x2_0_Output_01.write
		.adaptor_2x2_0_Output_01_writedata               (mm_interconnect_1_adaptor_2x2_0_output_01_writedata),          //                                          .writedata
		.adaptor_2x2_0_Output_01_waitrequest             (mm_interconnect_1_adaptor_2x2_0_output_01_waitrequest),        //                                          .waitrequest
		.Data_Memory_01_s1_address                       (mm_interconnect_1_data_memory_01_s1_address),                  //                         Data_Memory_01_s1.address
		.Data_Memory_01_s1_write                         (mm_interconnect_1_data_memory_01_s1_write),                    //                                          .write
		.Data_Memory_01_s1_readdata                      (mm_interconnect_1_data_memory_01_s1_readdata),                 //                                          .readdata
		.Data_Memory_01_s1_writedata                     (mm_interconnect_1_data_memory_01_s1_writedata),                //                                          .writedata
		.Data_Memory_01_s1_byteenable                    (mm_interconnect_1_data_memory_01_s1_byteenable),               //                                          .byteenable
		.Data_Memory_01_s1_chipselect                    (mm_interconnect_1_data_memory_01_s1_chipselect),               //                                          .chipselect
		.Data_Memory_01_s1_clken                         (mm_interconnect_1_data_memory_01_s1_clken),                    //                                          .clken
		.Instruction_Memory_01_s1_address                (mm_interconnect_1_instruction_memory_01_s1_address),           //                  Instruction_Memory_01_s1.address
		.Instruction_Memory_01_s1_write                  (mm_interconnect_1_instruction_memory_01_s1_write),             //                                          .write
		.Instruction_Memory_01_s1_readdata               (mm_interconnect_1_instruction_memory_01_s1_readdata),          //                                          .readdata
		.Instruction_Memory_01_s1_writedata              (mm_interconnect_1_instruction_memory_01_s1_writedata),         //                                          .writedata
		.Instruction_Memory_01_s1_byteenable             (mm_interconnect_1_instruction_memory_01_s1_byteenable),        //                                          .byteenable
		.Instruction_Memory_01_s1_chipselect             (mm_interconnect_1_instruction_memory_01_s1_chipselect),        //                                          .chipselect
		.Instruction_Memory_01_s1_clken                  (mm_interconnect_1_instruction_memory_01_s1_clken),             //                                          .clken
		.jtag_uart_01_avalon_jtag_slave_address          (mm_interconnect_1_jtag_uart_01_avalon_jtag_slave_address),     //            jtag_uart_01_avalon_jtag_slave.address
		.jtag_uart_01_avalon_jtag_slave_write            (mm_interconnect_1_jtag_uart_01_avalon_jtag_slave_write),       //                                          .write
		.jtag_uart_01_avalon_jtag_slave_read             (mm_interconnect_1_jtag_uart_01_avalon_jtag_slave_read),        //                                          .read
		.jtag_uart_01_avalon_jtag_slave_readdata         (mm_interconnect_1_jtag_uart_01_avalon_jtag_slave_readdata),    //                                          .readdata
		.jtag_uart_01_avalon_jtag_slave_writedata        (mm_interconnect_1_jtag_uart_01_avalon_jtag_slave_writedata),   //                                          .writedata
		.jtag_uart_01_avalon_jtag_slave_waitrequest      (mm_interconnect_1_jtag_uart_01_avalon_jtag_slave_waitrequest), //                                          .waitrequest
		.jtag_uart_01_avalon_jtag_slave_chipselect       (mm_interconnect_1_jtag_uart_01_avalon_jtag_slave_chipselect),  //                                          .chipselect
		.nios2_gen2_01_debug_mem_slave_address           (mm_interconnect_1_nios2_gen2_01_debug_mem_slave_address),      //             nios2_gen2_01_debug_mem_slave.address
		.nios2_gen2_01_debug_mem_slave_write             (mm_interconnect_1_nios2_gen2_01_debug_mem_slave_write),        //                                          .write
		.nios2_gen2_01_debug_mem_slave_read              (mm_interconnect_1_nios2_gen2_01_debug_mem_slave_read),         //                                          .read
		.nios2_gen2_01_debug_mem_slave_readdata          (mm_interconnect_1_nios2_gen2_01_debug_mem_slave_readdata),     //                                          .readdata
		.nios2_gen2_01_debug_mem_slave_writedata         (mm_interconnect_1_nios2_gen2_01_debug_mem_slave_writedata),    //                                          .writedata
		.nios2_gen2_01_debug_mem_slave_byteenable        (mm_interconnect_1_nios2_gen2_01_debug_mem_slave_byteenable),   //                                          .byteenable
		.nios2_gen2_01_debug_mem_slave_waitrequest       (mm_interconnect_1_nios2_gen2_01_debug_mem_slave_waitrequest),  //                                          .waitrequest
		.nios2_gen2_01_debug_mem_slave_debugaccess       (mm_interconnect_1_nios2_gen2_01_debug_mem_slave_debugaccess)   //                                          .debugaccess
	);

	adaptor2x2_mm_interconnect_2 mm_interconnect_2 (
		.clk_0_clk_clk                                   (clk_clk),                                                      //                                 clk_0_clk.clk
		.nios2_gen2_10_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                               // nios2_gen2_10_reset_reset_bridge_in_reset.reset
		.nios2_gen2_10_data_master_address               (nios2_gen2_10_data_master_address),                            //                 nios2_gen2_10_data_master.address
		.nios2_gen2_10_data_master_waitrequest           (nios2_gen2_10_data_master_waitrequest),                        //                                          .waitrequest
		.nios2_gen2_10_data_master_byteenable            (nios2_gen2_10_data_master_byteenable),                         //                                          .byteenable
		.nios2_gen2_10_data_master_read                  (nios2_gen2_10_data_master_read),                               //                                          .read
		.nios2_gen2_10_data_master_readdata              (nios2_gen2_10_data_master_readdata),                           //                                          .readdata
		.nios2_gen2_10_data_master_write                 (nios2_gen2_10_data_master_write),                              //                                          .write
		.nios2_gen2_10_data_master_writedata             (nios2_gen2_10_data_master_writedata),                          //                                          .writedata
		.nios2_gen2_10_data_master_debugaccess           (nios2_gen2_10_data_master_debugaccess),                        //                                          .debugaccess
		.nios2_gen2_10_instruction_master_address        (nios2_gen2_10_instruction_master_address),                     //          nios2_gen2_10_instruction_master.address
		.nios2_gen2_10_instruction_master_waitrequest    (nios2_gen2_10_instruction_master_waitrequest),                 //                                          .waitrequest
		.nios2_gen2_10_instruction_master_read           (nios2_gen2_10_instruction_master_read),                        //                                          .read
		.nios2_gen2_10_instruction_master_readdata       (nios2_gen2_10_instruction_master_readdata),                    //                                          .readdata
		.adaptor_2x2_0_Input_10_read                     (mm_interconnect_2_adaptor_2x2_0_input_10_read),                //                    adaptor_2x2_0_Input_10.read
		.adaptor_2x2_0_Input_10_readdata                 (mm_interconnect_2_adaptor_2x2_0_input_10_readdata),            //                                          .readdata
		.adaptor_2x2_0_Output_10_write                   (mm_interconnect_2_adaptor_2x2_0_output_10_write),              //                   adaptor_2x2_0_Output_10.write
		.adaptor_2x2_0_Output_10_writedata               (mm_interconnect_2_adaptor_2x2_0_output_10_writedata),          //                                          .writedata
		.adaptor_2x2_0_Output_10_waitrequest             (mm_interconnect_2_adaptor_2x2_0_output_10_waitrequest),        //                                          .waitrequest
		.Data_Memory_10_s1_address                       (mm_interconnect_2_data_memory_10_s1_address),                  //                         Data_Memory_10_s1.address
		.Data_Memory_10_s1_write                         (mm_interconnect_2_data_memory_10_s1_write),                    //                                          .write
		.Data_Memory_10_s1_readdata                      (mm_interconnect_2_data_memory_10_s1_readdata),                 //                                          .readdata
		.Data_Memory_10_s1_writedata                     (mm_interconnect_2_data_memory_10_s1_writedata),                //                                          .writedata
		.Data_Memory_10_s1_byteenable                    (mm_interconnect_2_data_memory_10_s1_byteenable),               //                                          .byteenable
		.Data_Memory_10_s1_chipselect                    (mm_interconnect_2_data_memory_10_s1_chipselect),               //                                          .chipselect
		.Data_Memory_10_s1_clken                         (mm_interconnect_2_data_memory_10_s1_clken),                    //                                          .clken
		.Instruction_Memory_10_s1_address                (mm_interconnect_2_instruction_memory_10_s1_address),           //                  Instruction_Memory_10_s1.address
		.Instruction_Memory_10_s1_write                  (mm_interconnect_2_instruction_memory_10_s1_write),             //                                          .write
		.Instruction_Memory_10_s1_readdata               (mm_interconnect_2_instruction_memory_10_s1_readdata),          //                                          .readdata
		.Instruction_Memory_10_s1_writedata              (mm_interconnect_2_instruction_memory_10_s1_writedata),         //                                          .writedata
		.Instruction_Memory_10_s1_byteenable             (mm_interconnect_2_instruction_memory_10_s1_byteenable),        //                                          .byteenable
		.Instruction_Memory_10_s1_chipselect             (mm_interconnect_2_instruction_memory_10_s1_chipselect),        //                                          .chipselect
		.Instruction_Memory_10_s1_clken                  (mm_interconnect_2_instruction_memory_10_s1_clken),             //                                          .clken
		.jtag_uart_10_avalon_jtag_slave_address          (mm_interconnect_2_jtag_uart_10_avalon_jtag_slave_address),     //            jtag_uart_10_avalon_jtag_slave.address
		.jtag_uart_10_avalon_jtag_slave_write            (mm_interconnect_2_jtag_uart_10_avalon_jtag_slave_write),       //                                          .write
		.jtag_uart_10_avalon_jtag_slave_read             (mm_interconnect_2_jtag_uart_10_avalon_jtag_slave_read),        //                                          .read
		.jtag_uart_10_avalon_jtag_slave_readdata         (mm_interconnect_2_jtag_uart_10_avalon_jtag_slave_readdata),    //                                          .readdata
		.jtag_uart_10_avalon_jtag_slave_writedata        (mm_interconnect_2_jtag_uart_10_avalon_jtag_slave_writedata),   //                                          .writedata
		.jtag_uart_10_avalon_jtag_slave_waitrequest      (mm_interconnect_2_jtag_uart_10_avalon_jtag_slave_waitrequest), //                                          .waitrequest
		.jtag_uart_10_avalon_jtag_slave_chipselect       (mm_interconnect_2_jtag_uart_10_avalon_jtag_slave_chipselect),  //                                          .chipselect
		.nios2_gen2_10_debug_mem_slave_address           (mm_interconnect_2_nios2_gen2_10_debug_mem_slave_address),      //             nios2_gen2_10_debug_mem_slave.address
		.nios2_gen2_10_debug_mem_slave_write             (mm_interconnect_2_nios2_gen2_10_debug_mem_slave_write),        //                                          .write
		.nios2_gen2_10_debug_mem_slave_read              (mm_interconnect_2_nios2_gen2_10_debug_mem_slave_read),         //                                          .read
		.nios2_gen2_10_debug_mem_slave_readdata          (mm_interconnect_2_nios2_gen2_10_debug_mem_slave_readdata),     //                                          .readdata
		.nios2_gen2_10_debug_mem_slave_writedata         (mm_interconnect_2_nios2_gen2_10_debug_mem_slave_writedata),    //                                          .writedata
		.nios2_gen2_10_debug_mem_slave_byteenable        (mm_interconnect_2_nios2_gen2_10_debug_mem_slave_byteenable),   //                                          .byteenable
		.nios2_gen2_10_debug_mem_slave_waitrequest       (mm_interconnect_2_nios2_gen2_10_debug_mem_slave_waitrequest),  //                                          .waitrequest
		.nios2_gen2_10_debug_mem_slave_debugaccess       (mm_interconnect_2_nios2_gen2_10_debug_mem_slave_debugaccess)   //                                          .debugaccess
	);

	adaptor2x2_mm_interconnect_3 mm_interconnect_3 (
		.clk_0_clk_clk                                   (clk_clk),                                                      //                                 clk_0_clk.clk
		.nios2_gen2_11_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                               // nios2_gen2_11_reset_reset_bridge_in_reset.reset
		.nios2_gen2_11_data_master_address               (nios2_gen2_11_data_master_address),                            //                 nios2_gen2_11_data_master.address
		.nios2_gen2_11_data_master_waitrequest           (nios2_gen2_11_data_master_waitrequest),                        //                                          .waitrequest
		.nios2_gen2_11_data_master_byteenable            (nios2_gen2_11_data_master_byteenable),                         //                                          .byteenable
		.nios2_gen2_11_data_master_read                  (nios2_gen2_11_data_master_read),                               //                                          .read
		.nios2_gen2_11_data_master_readdata              (nios2_gen2_11_data_master_readdata),                           //                                          .readdata
		.nios2_gen2_11_data_master_write                 (nios2_gen2_11_data_master_write),                              //                                          .write
		.nios2_gen2_11_data_master_writedata             (nios2_gen2_11_data_master_writedata),                          //                                          .writedata
		.nios2_gen2_11_data_master_debugaccess           (nios2_gen2_11_data_master_debugaccess),                        //                                          .debugaccess
		.nios2_gen2_11_instruction_master_address        (nios2_gen2_11_instruction_master_address),                     //          nios2_gen2_11_instruction_master.address
		.nios2_gen2_11_instruction_master_waitrequest    (nios2_gen2_11_instruction_master_waitrequest),                 //                                          .waitrequest
		.nios2_gen2_11_instruction_master_read           (nios2_gen2_11_instruction_master_read),                        //                                          .read
		.nios2_gen2_11_instruction_master_readdata       (nios2_gen2_11_instruction_master_readdata),                    //                                          .readdata
		.adaptor_2x2_0_Input_11_read                     (mm_interconnect_3_adaptor_2x2_0_input_11_read),                //                    adaptor_2x2_0_Input_11.read
		.adaptor_2x2_0_Input_11_readdata                 (mm_interconnect_3_adaptor_2x2_0_input_11_readdata),            //                                          .readdata
		.adaptor_2x2_0_Output_11_write                   (mm_interconnect_3_adaptor_2x2_0_output_11_write),              //                   adaptor_2x2_0_Output_11.write
		.adaptor_2x2_0_Output_11_writedata               (mm_interconnect_3_adaptor_2x2_0_output_11_writedata),          //                                          .writedata
		.adaptor_2x2_0_Output_11_waitrequest             (mm_interconnect_3_adaptor_2x2_0_output_11_waitrequest),        //                                          .waitrequest
		.Data_Memory_11_s1_address                       (mm_interconnect_3_data_memory_11_s1_address),                  //                         Data_Memory_11_s1.address
		.Data_Memory_11_s1_write                         (mm_interconnect_3_data_memory_11_s1_write),                    //                                          .write
		.Data_Memory_11_s1_readdata                      (mm_interconnect_3_data_memory_11_s1_readdata),                 //                                          .readdata
		.Data_Memory_11_s1_writedata                     (mm_interconnect_3_data_memory_11_s1_writedata),                //                                          .writedata
		.Data_Memory_11_s1_byteenable                    (mm_interconnect_3_data_memory_11_s1_byteenable),               //                                          .byteenable
		.Data_Memory_11_s1_chipselect                    (mm_interconnect_3_data_memory_11_s1_chipselect),               //                                          .chipselect
		.Data_Memory_11_s1_clken                         (mm_interconnect_3_data_memory_11_s1_clken),                    //                                          .clken
		.Instruction_Memory_11_s1_address                (mm_interconnect_3_instruction_memory_11_s1_address),           //                  Instruction_Memory_11_s1.address
		.Instruction_Memory_11_s1_write                  (mm_interconnect_3_instruction_memory_11_s1_write),             //                                          .write
		.Instruction_Memory_11_s1_readdata               (mm_interconnect_3_instruction_memory_11_s1_readdata),          //                                          .readdata
		.Instruction_Memory_11_s1_writedata              (mm_interconnect_3_instruction_memory_11_s1_writedata),         //                                          .writedata
		.Instruction_Memory_11_s1_byteenable             (mm_interconnect_3_instruction_memory_11_s1_byteenable),        //                                          .byteenable
		.Instruction_Memory_11_s1_chipselect             (mm_interconnect_3_instruction_memory_11_s1_chipselect),        //                                          .chipselect
		.Instruction_Memory_11_s1_clken                  (mm_interconnect_3_instruction_memory_11_s1_clken),             //                                          .clken
		.jtag_uart_11_avalon_jtag_slave_address          (mm_interconnect_3_jtag_uart_11_avalon_jtag_slave_address),     //            jtag_uart_11_avalon_jtag_slave.address
		.jtag_uart_11_avalon_jtag_slave_write            (mm_interconnect_3_jtag_uart_11_avalon_jtag_slave_write),       //                                          .write
		.jtag_uart_11_avalon_jtag_slave_read             (mm_interconnect_3_jtag_uart_11_avalon_jtag_slave_read),        //                                          .read
		.jtag_uart_11_avalon_jtag_slave_readdata         (mm_interconnect_3_jtag_uart_11_avalon_jtag_slave_readdata),    //                                          .readdata
		.jtag_uart_11_avalon_jtag_slave_writedata        (mm_interconnect_3_jtag_uart_11_avalon_jtag_slave_writedata),   //                                          .writedata
		.jtag_uart_11_avalon_jtag_slave_waitrequest      (mm_interconnect_3_jtag_uart_11_avalon_jtag_slave_waitrequest), //                                          .waitrequest
		.jtag_uart_11_avalon_jtag_slave_chipselect       (mm_interconnect_3_jtag_uart_11_avalon_jtag_slave_chipselect),  //                                          .chipselect
		.nios2_gen2_11_debug_mem_slave_address           (mm_interconnect_3_nios2_gen2_11_debug_mem_slave_address),      //             nios2_gen2_11_debug_mem_slave.address
		.nios2_gen2_11_debug_mem_slave_write             (mm_interconnect_3_nios2_gen2_11_debug_mem_slave_write),        //                                          .write
		.nios2_gen2_11_debug_mem_slave_read              (mm_interconnect_3_nios2_gen2_11_debug_mem_slave_read),         //                                          .read
		.nios2_gen2_11_debug_mem_slave_readdata          (mm_interconnect_3_nios2_gen2_11_debug_mem_slave_readdata),     //                                          .readdata
		.nios2_gen2_11_debug_mem_slave_writedata         (mm_interconnect_3_nios2_gen2_11_debug_mem_slave_writedata),    //                                          .writedata
		.nios2_gen2_11_debug_mem_slave_byteenable        (mm_interconnect_3_nios2_gen2_11_debug_mem_slave_byteenable),   //                                          .byteenable
		.nios2_gen2_11_debug_mem_slave_waitrequest       (mm_interconnect_3_nios2_gen2_11_debug_mem_slave_waitrequest),  //                                          .waitrequest
		.nios2_gen2_11_debug_mem_slave_debugaccess       (mm_interconnect_3_nios2_gen2_11_debug_mem_slave_debugaccess)   //                                          .debugaccess
	);

	adaptor2x2_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (nios2_gen2_00_irq_irq)           //    sender.irq
	);

	adaptor2x2_irq_mapper irq_mapper_001 (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_001_receiver0_irq),   // receiver0.irq
		.receiver1_irq (irq_mapper_001_receiver1_irq),   // receiver1.irq
		.sender_irq    (nios2_gen2_01_irq_irq)           //    sender.irq
	);

	adaptor2x2_irq_mapper irq_mapper_002 (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_002_receiver0_irq),   // receiver0.irq
		.receiver1_irq (irq_mapper_002_receiver1_irq),   // receiver1.irq
		.sender_irq    (nios2_gen2_10_irq_irq)           //    sender.irq
	);

	adaptor2x2_irq_mapper irq_mapper_003 (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_003_receiver0_irq),   // receiver0.irq
		.receiver1_irq (irq_mapper_003_receiver1_irq),   // receiver1.irq
		.sender_irq    (nios2_gen2_11_irq_irq)           //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
