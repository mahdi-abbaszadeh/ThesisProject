
module NoC_QSYS (
	clk_clk);	

	input		clk_clk;
endmodule
