
module adaptor2x2 (
	reset_reset_n,
	clk_clk);	

	input		reset_reset_n;
	input		clk_clk;
endmodule
