// unsaved.v

// Generated using ACDS version 17.1 590

`timescale 1 ps / 1 ps
module unsaved (
		input  wire  clk_clk,       //   clk.clk
		input  wire  reset_reset_n  // reset.reset_n
	);

	wire         mm2stfifo_0_out_valid;                                       // MM2STFIFO_0:avalonst_source_valid -> ST2MMFIFO_1:avalonst_sink_valid
	wire  [31:0] mm2stfifo_0_out_data;                                        // MM2STFIFO_0:avalonst_source_data -> ST2MMFIFO_1:avalonst_sink_data
	wire         mm2stfifo_0_out_ready;                                       // ST2MMFIFO_1:avalonst_sink_ready -> MM2STFIFO_0:avalonst_source_ready
	wire   [7:0] mm2stfifo_0_out_channel;                                     // MM2STFIFO_0:avalonst_source_channel -> ST2MMFIFO_1:avalonst_sink_channel
	wire   [7:0] mm2stfifo_0_out_error;                                       // MM2STFIFO_0:avalonst_source_error -> ST2MMFIFO_1:avalonst_sink_error
	wire         mm2stfifo_1_out_valid;                                       // MM2STFIFO_1:avalonst_source_valid -> ST2MMFIFO_0:avalonst_sink_valid
	wire  [31:0] mm2stfifo_1_out_data;                                        // MM2STFIFO_1:avalonst_source_data -> ST2MMFIFO_0:avalonst_sink_data
	wire         mm2stfifo_1_out_ready;                                       // ST2MMFIFO_0:avalonst_sink_ready -> MM2STFIFO_1:avalonst_source_ready
	wire   [7:0] mm2stfifo_1_out_channel;                                     // MM2STFIFO_1:avalonst_source_channel -> ST2MMFIFO_0:avalonst_sink_channel
	wire   [7:0] mm2stfifo_1_out_error;                                       // MM2STFIFO_1:avalonst_source_error -> ST2MMFIFO_0:avalonst_sink_error
	wire  [31:0] nios2_gen2_0_data_master_readdata;                           // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                        // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                        // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [17:0] nios2_gen2_0_data_master_address;                            // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                         // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                               // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_write;                              // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                          // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire  [31:0] nios2_gen2_1_data_master_readdata;                           // mm_interconnect_0:nios2_gen2_1_data_master_readdata -> nios2_gen2_1:d_readdata
	wire         nios2_gen2_1_data_master_waitrequest;                        // mm_interconnect_0:nios2_gen2_1_data_master_waitrequest -> nios2_gen2_1:d_waitrequest
	wire         nios2_gen2_1_data_master_debugaccess;                        // nios2_gen2_1:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_1_data_master_debugaccess
	wire  [17:0] nios2_gen2_1_data_master_address;                            // nios2_gen2_1:d_address -> mm_interconnect_0:nios2_gen2_1_data_master_address
	wire   [3:0] nios2_gen2_1_data_master_byteenable;                         // nios2_gen2_1:d_byteenable -> mm_interconnect_0:nios2_gen2_1_data_master_byteenable
	wire         nios2_gen2_1_data_master_read;                               // nios2_gen2_1:d_read -> mm_interconnect_0:nios2_gen2_1_data_master_read
	wire         nios2_gen2_1_data_master_write;                              // nios2_gen2_1:d_write -> mm_interconnect_0:nios2_gen2_1_data_master_write
	wire  [31:0] nios2_gen2_1_data_master_writedata;                          // nios2_gen2_1:d_writedata -> mm_interconnect_0:nios2_gen2_1_data_master_writedata
	wire  [31:0] nios2_gen2_1_instruction_master_readdata;                    // mm_interconnect_0:nios2_gen2_1_instruction_master_readdata -> nios2_gen2_1:i_readdata
	wire         nios2_gen2_1_instruction_master_waitrequest;                 // mm_interconnect_0:nios2_gen2_1_instruction_master_waitrequest -> nios2_gen2_1:i_waitrequest
	wire  [17:0] nios2_gen2_1_instruction_master_address;                     // nios2_gen2_1:i_address -> mm_interconnect_0:nios2_gen2_1_instruction_master_address
	wire         nios2_gen2_1_instruction_master_read;                        // nios2_gen2_1:i_read -> mm_interconnect_0:nios2_gen2_1_instruction_master_read
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                    // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                 // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [17:0] nios2_gen2_0_instruction_master_address;                     // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                        // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;     // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest;  // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess;  // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;      // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;         // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;   // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;        // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;    // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire         mm_interconnect_0_mm2stfifo_0_in_waitrequest;                // MM2STFIFO_0:avalonmm_write_slave_waitrequest -> mm_interconnect_0:MM2STFIFO_0_in_waitrequest
	wire   [0:0] mm_interconnect_0_mm2stfifo_0_in_address;                    // mm_interconnect_0:MM2STFIFO_0_in_address -> MM2STFIFO_0:avalonmm_write_slave_address
	wire         mm_interconnect_0_mm2stfifo_0_in_write;                      // mm_interconnect_0:MM2STFIFO_0_in_write -> MM2STFIFO_0:avalonmm_write_slave_write
	wire  [31:0] mm_interconnect_0_mm2stfifo_0_in_writedata;                  // mm_interconnect_0:MM2STFIFO_0_in_writedata -> MM2STFIFO_0:avalonmm_write_slave_writedata
	wire  [31:0] mm_interconnect_0_mm2stfifo_0_in_csr_readdata;               // MM2STFIFO_0:wrclk_control_slave_readdata -> mm_interconnect_0:MM2STFIFO_0_in_csr_readdata
	wire   [2:0] mm_interconnect_0_mm2stfifo_0_in_csr_address;                // mm_interconnect_0:MM2STFIFO_0_in_csr_address -> MM2STFIFO_0:wrclk_control_slave_address
	wire         mm_interconnect_0_mm2stfifo_0_in_csr_read;                   // mm_interconnect_0:MM2STFIFO_0_in_csr_read -> MM2STFIFO_0:wrclk_control_slave_read
	wire         mm_interconnect_0_mm2stfifo_0_in_csr_write;                  // mm_interconnect_0:MM2STFIFO_0_in_csr_write -> MM2STFIFO_0:wrclk_control_slave_write
	wire  [31:0] mm_interconnect_0_mm2stfifo_0_in_csr_writedata;              // mm_interconnect_0:MM2STFIFO_0_in_csr_writedata -> MM2STFIFO_0:wrclk_control_slave_writedata
	wire  [31:0] mm_interconnect_0_st2mmfifo_0_in_csr_readdata;               // ST2MMFIFO_0:wrclk_control_slave_readdata -> mm_interconnect_0:ST2MMFIFO_0_in_csr_readdata
	wire   [2:0] mm_interconnect_0_st2mmfifo_0_in_csr_address;                // mm_interconnect_0:ST2MMFIFO_0_in_csr_address -> ST2MMFIFO_0:wrclk_control_slave_address
	wire         mm_interconnect_0_st2mmfifo_0_in_csr_read;                   // mm_interconnect_0:ST2MMFIFO_0_in_csr_read -> ST2MMFIFO_0:wrclk_control_slave_read
	wire         mm_interconnect_0_st2mmfifo_0_in_csr_write;                  // mm_interconnect_0:ST2MMFIFO_0_in_csr_write -> ST2MMFIFO_0:wrclk_control_slave_write
	wire  [31:0] mm_interconnect_0_st2mmfifo_0_in_csr_writedata;              // mm_interconnect_0:ST2MMFIFO_0_in_csr_writedata -> ST2MMFIFO_0:wrclk_control_slave_writedata
	wire  [31:0] mm_interconnect_0_st2mmfifo_0_out_readdata;                  // ST2MMFIFO_0:avalonmm_read_slave_readdata -> mm_interconnect_0:ST2MMFIFO_0_out_readdata
	wire         mm_interconnect_0_st2mmfifo_0_out_waitrequest;               // ST2MMFIFO_0:avalonmm_read_slave_waitrequest -> mm_interconnect_0:ST2MMFIFO_0_out_waitrequest
	wire   [0:0] mm_interconnect_0_st2mmfifo_0_out_address;                   // mm_interconnect_0:ST2MMFIFO_0_out_address -> ST2MMFIFO_0:avalonmm_read_slave_address
	wire         mm_interconnect_0_st2mmfifo_0_out_read;                      // mm_interconnect_0:ST2MMFIFO_0_out_read -> ST2MMFIFO_0:avalonmm_read_slave_read
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;            // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;              // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire  [13:0] mm_interconnect_0_onchip_memory2_0_s1_address;               // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;            // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                 // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;             // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                 // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire  [31:0] mm_interconnect_0_nios2_gen2_1_debug_mem_slave_readdata;     // nios2_gen2_1:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_1_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_1_debug_mem_slave_waitrequest;  // nios2_gen2_1:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_1_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_1_debug_mem_slave_debugaccess;  // mm_interconnect_0:nios2_gen2_1_debug_mem_slave_debugaccess -> nios2_gen2_1:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_1_debug_mem_slave_address;      // mm_interconnect_0:nios2_gen2_1_debug_mem_slave_address -> nios2_gen2_1:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_1_debug_mem_slave_read;         // mm_interconnect_0:nios2_gen2_1_debug_mem_slave_read -> nios2_gen2_1:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_1_debug_mem_slave_byteenable;   // mm_interconnect_0:nios2_gen2_1_debug_mem_slave_byteenable -> nios2_gen2_1:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_1_debug_mem_slave_write;        // mm_interconnect_0:nios2_gen2_1_debug_mem_slave_write -> nios2_gen2_1:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_1_debug_mem_slave_writedata;    // mm_interconnect_0:nios2_gen2_1_debug_mem_slave_writedata -> nios2_gen2_1:debug_mem_slave_writedata
	wire         mm_interconnect_0_mm2stfifo_1_in_waitrequest;                // MM2STFIFO_1:avalonmm_write_slave_waitrequest -> mm_interconnect_0:MM2STFIFO_1_in_waitrequest
	wire   [0:0] mm_interconnect_0_mm2stfifo_1_in_address;                    // mm_interconnect_0:MM2STFIFO_1_in_address -> MM2STFIFO_1:avalonmm_write_slave_address
	wire         mm_interconnect_0_mm2stfifo_1_in_write;                      // mm_interconnect_0:MM2STFIFO_1_in_write -> MM2STFIFO_1:avalonmm_write_slave_write
	wire  [31:0] mm_interconnect_0_mm2stfifo_1_in_writedata;                  // mm_interconnect_0:MM2STFIFO_1_in_writedata -> MM2STFIFO_1:avalonmm_write_slave_writedata
	wire  [31:0] mm_interconnect_0_st2mmfifo_1_in_csr_readdata;               // ST2MMFIFO_1:wrclk_control_slave_readdata -> mm_interconnect_0:ST2MMFIFO_1_in_csr_readdata
	wire   [2:0] mm_interconnect_0_st2mmfifo_1_in_csr_address;                // mm_interconnect_0:ST2MMFIFO_1_in_csr_address -> ST2MMFIFO_1:wrclk_control_slave_address
	wire         mm_interconnect_0_st2mmfifo_1_in_csr_read;                   // mm_interconnect_0:ST2MMFIFO_1_in_csr_read -> ST2MMFIFO_1:wrclk_control_slave_read
	wire         mm_interconnect_0_st2mmfifo_1_in_csr_write;                  // mm_interconnect_0:ST2MMFIFO_1_in_csr_write -> ST2MMFIFO_1:wrclk_control_slave_write
	wire  [31:0] mm_interconnect_0_st2mmfifo_1_in_csr_writedata;              // mm_interconnect_0:ST2MMFIFO_1_in_csr_writedata -> ST2MMFIFO_1:wrclk_control_slave_writedata
	wire  [31:0] mm_interconnect_0_mm2stfifo_1_in_csr_readdata;               // MM2STFIFO_1:wrclk_control_slave_readdata -> mm_interconnect_0:MM2STFIFO_1_in_csr_readdata
	wire   [2:0] mm_interconnect_0_mm2stfifo_1_in_csr_address;                // mm_interconnect_0:MM2STFIFO_1_in_csr_address -> MM2STFIFO_1:wrclk_control_slave_address
	wire         mm_interconnect_0_mm2stfifo_1_in_csr_read;                   // mm_interconnect_0:MM2STFIFO_1_in_csr_read -> MM2STFIFO_1:wrclk_control_slave_read
	wire         mm_interconnect_0_mm2stfifo_1_in_csr_write;                  // mm_interconnect_0:MM2STFIFO_1_in_csr_write -> MM2STFIFO_1:wrclk_control_slave_write
	wire  [31:0] mm_interconnect_0_mm2stfifo_1_in_csr_writedata;              // mm_interconnect_0:MM2STFIFO_1_in_csr_writedata -> MM2STFIFO_1:wrclk_control_slave_writedata
	wire  [31:0] mm_interconnect_0_st2mmfifo_1_out_readdata;                  // ST2MMFIFO_1:avalonmm_read_slave_readdata -> mm_interconnect_0:ST2MMFIFO_1_out_readdata
	wire         mm_interconnect_0_st2mmfifo_1_out_waitrequest;               // ST2MMFIFO_1:avalonmm_read_slave_waitrequest -> mm_interconnect_0:ST2MMFIFO_1_out_waitrequest
	wire   [0:0] mm_interconnect_0_st2mmfifo_1_out_address;                   // mm_interconnect_0:ST2MMFIFO_1_out_address -> ST2MMFIFO_1:avalonmm_read_slave_address
	wire         mm_interconnect_0_st2mmfifo_1_out_read;                      // mm_interconnect_0:ST2MMFIFO_1_out_read -> ST2MMFIFO_1:avalonmm_read_slave_read
	wire         mm_interconnect_0_onchip_memory2_1_s1_chipselect;            // mm_interconnect_0:onchip_memory2_1_s1_chipselect -> onchip_memory2_1:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_1_s1_readdata;              // onchip_memory2_1:readdata -> mm_interconnect_0:onchip_memory2_1_s1_readdata
	wire  [13:0] mm_interconnect_0_onchip_memory2_1_s1_address;               // mm_interconnect_0:onchip_memory2_1_s1_address -> onchip_memory2_1:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_1_s1_byteenable;            // mm_interconnect_0:onchip_memory2_1_s1_byteenable -> onchip_memory2_1:byteenable
	wire         mm_interconnect_0_onchip_memory2_1_s1_write;                 // mm_interconnect_0:onchip_memory2_1_s1_write -> onchip_memory2_1:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_1_s1_writedata;             // mm_interconnect_0:onchip_memory2_1_s1_writedata -> onchip_memory2_1:writedata
	wire         mm_interconnect_0_onchip_memory2_1_s1_clken;                 // mm_interconnect_0:onchip_memory2_1_s1_clken -> onchip_memory2_1:clken
	wire         mm_interconnect_0_inst_mem_1_s1_chipselect;                  // mm_interconnect_0:Inst_mem_1_s1_chipselect -> Inst_mem_1:chipselect
	wire  [31:0] mm_interconnect_0_inst_mem_1_s1_readdata;                    // Inst_mem_1:readdata -> mm_interconnect_0:Inst_mem_1_s1_readdata
	wire  [13:0] mm_interconnect_0_inst_mem_1_s1_address;                     // mm_interconnect_0:Inst_mem_1_s1_address -> Inst_mem_1:address
	wire   [3:0] mm_interconnect_0_inst_mem_1_s1_byteenable;                  // mm_interconnect_0:Inst_mem_1_s1_byteenable -> Inst_mem_1:byteenable
	wire         mm_interconnect_0_inst_mem_1_s1_write;                       // mm_interconnect_0:Inst_mem_1_s1_write -> Inst_mem_1:write
	wire  [31:0] mm_interconnect_0_inst_mem_1_s1_writedata;                   // mm_interconnect_0:Inst_mem_1_s1_writedata -> Inst_mem_1:writedata
	wire         mm_interconnect_0_inst_mem_1_s1_clken;                       // mm_interconnect_0:Inst_mem_1_s1_clken -> Inst_mem_1:clken
	wire         mm_interconnect_0_inst_mem_0_s1_chipselect;                  // mm_interconnect_0:Inst_mem_0_s1_chipselect -> Inst_mem_0:chipselect
	wire  [31:0] mm_interconnect_0_inst_mem_0_s1_readdata;                    // Inst_mem_0:readdata -> mm_interconnect_0:Inst_mem_0_s1_readdata
	wire  [13:0] mm_interconnect_0_inst_mem_0_s1_address;                     // mm_interconnect_0:Inst_mem_0_s1_address -> Inst_mem_0:address
	wire   [3:0] mm_interconnect_0_inst_mem_0_s1_byteenable;                  // mm_interconnect_0:Inst_mem_0_s1_byteenable -> Inst_mem_0:byteenable
	wire         mm_interconnect_0_inst_mem_0_s1_write;                       // mm_interconnect_0:Inst_mem_0_s1_write -> Inst_mem_0:write
	wire  [31:0] mm_interconnect_0_inst_mem_0_s1_writedata;                   // mm_interconnect_0:Inst_mem_0_s1_writedata -> Inst_mem_0:writedata
	wire         mm_interconnect_0_inst_mem_0_s1_clken;                       // mm_interconnect_0:Inst_mem_0_s1_clken -> Inst_mem_0:clken
	wire         irq_mapper_receiver0_irq;                                    // MM2STFIFO_0:wrclk_control_slave_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                    // ST2MMFIFO_0:wrclk_control_slave_irq -> irq_mapper:receiver1_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                        // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         irq_mapper_001_receiver0_irq;                                // MM2STFIFO_1:wrclk_control_slave_irq -> irq_mapper_001:receiver0_irq
	wire         irq_mapper_001_receiver1_irq;                                // ST2MMFIFO_1:wrclk_control_slave_irq -> irq_mapper_001:receiver1_irq
	wire  [31:0] nios2_gen2_1_irq_irq;                                        // irq_mapper_001:sender_irq -> nios2_gen2_1:irq
	wire         irq_mapper_receiver2_irq;                                    // jtag_uart_0:av_irq -> [irq_mapper:receiver2_irq, irq_mapper_001:receiver2_irq]
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [Inst_mem_0:reset, Inst_mem_1:reset, MM2STFIFO_0:reset_n, MM2STFIFO_1:reset_n, ST2MMFIFO_0:reset_n, ST2MMFIFO_1:reset_n, irq_mapper:reset, irq_mapper_001:reset, jtag_uart_0:rst_n, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n, nios2_gen2_1:reset_n, onchip_memory2_0:reset, onchip_memory2_1:reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                          // rst_controller:reset_req -> [Inst_mem_0:reset_req, Inst_mem_1:reset_req, nios2_gen2_0:reset_req, nios2_gen2_1:reset_req, onchip_memory2_0:reset_req, onchip_memory2_1:reset_req, rst_translator:reset_req_in]

	unsaved_Inst_mem_0 inst_mem_0 (
		.clk        (clk_clk),                                    //   clk1.clk
		.address    (mm_interconnect_0_inst_mem_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_inst_mem_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_inst_mem_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_inst_mem_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_inst_mem_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_inst_mem_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_inst_mem_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),             // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),         //       .reset_req
		.freeze     (1'b0)                                        // (terminated)
	);

	unsaved_Inst_mem_1 inst_mem_1 (
		.clk        (clk_clk),                                    //   clk1.clk
		.address    (mm_interconnect_0_inst_mem_1_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_inst_mem_1_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_inst_mem_1_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_inst_mem_1_s1_write),      //       .write
		.readdata   (mm_interconnect_0_inst_mem_1_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_inst_mem_1_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_inst_mem_1_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),             // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),         //       .reset_req
		.freeze     (1'b0)                                        // (terminated)
	);

	unsaved_MM2STFIFO_0 mm2stfifo_0 (
		.wrclock                          (clk_clk),                                        //   clk_in.clk
		.reset_n                          (~rst_controller_reset_out_reset),                // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_0_mm2stfifo_0_in_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_0_mm2stfifo_0_in_write),         //         .write
		.avalonmm_write_slave_address     (mm_interconnect_0_mm2stfifo_0_in_address),       //         .address
		.avalonmm_write_slave_waitrequest (mm_interconnect_0_mm2stfifo_0_in_waitrequest),   //         .waitrequest
		.avalonst_source_valid            (mm2stfifo_0_out_valid),                          //      out.valid
		.avalonst_source_data             (mm2stfifo_0_out_data),                           //         .data
		.avalonst_source_channel          (mm2stfifo_0_out_channel),                        //         .channel
		.avalonst_source_error            (mm2stfifo_0_out_error),                          //         .error
		.avalonst_source_ready            (mm2stfifo_0_out_ready),                          //         .ready
		.wrclk_control_slave_address      (mm_interconnect_0_mm2stfifo_0_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_0_mm2stfifo_0_in_csr_read),      //         .read
		.wrclk_control_slave_writedata    (mm_interconnect_0_mm2stfifo_0_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write        (mm_interconnect_0_mm2stfifo_0_in_csr_write),     //         .write
		.wrclk_control_slave_readdata     (mm_interconnect_0_mm2stfifo_0_in_csr_readdata),  //         .readdata
		.wrclk_control_slave_irq          (irq_mapper_receiver0_irq)                        //   in_irq.irq
	);

	unsaved_MM2STFIFO_0 mm2stfifo_1 (
		.wrclock                          (clk_clk),                                        //   clk_in.clk
		.reset_n                          (~rst_controller_reset_out_reset),                // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_0_mm2stfifo_1_in_writedata),     //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_0_mm2stfifo_1_in_write),         //         .write
		.avalonmm_write_slave_address     (mm_interconnect_0_mm2stfifo_1_in_address),       //         .address
		.avalonmm_write_slave_waitrequest (mm_interconnect_0_mm2stfifo_1_in_waitrequest),   //         .waitrequest
		.avalonst_source_valid            (mm2stfifo_1_out_valid),                          //      out.valid
		.avalonst_source_data             (mm2stfifo_1_out_data),                           //         .data
		.avalonst_source_channel          (mm2stfifo_1_out_channel),                        //         .channel
		.avalonst_source_error            (mm2stfifo_1_out_error),                          //         .error
		.avalonst_source_ready            (mm2stfifo_1_out_ready),                          //         .ready
		.wrclk_control_slave_address      (mm_interconnect_0_mm2stfifo_1_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read         (mm_interconnect_0_mm2stfifo_1_in_csr_read),      //         .read
		.wrclk_control_slave_writedata    (mm_interconnect_0_mm2stfifo_1_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write        (mm_interconnect_0_mm2stfifo_1_in_csr_write),     //         .write
		.wrclk_control_slave_readdata     (mm_interconnect_0_mm2stfifo_1_in_csr_readdata),  //         .readdata
		.wrclk_control_slave_irq          (irq_mapper_001_receiver0_irq)                    //   in_irq.irq
	);

	unsaved_ST2MMFIFO_0 st2mmfifo_0 (
		.wrclock                         (clk_clk),                                        //   clk_in.clk
		.reset_n                         (~rst_controller_reset_out_reset),                // reset_in.reset_n
		.avalonst_sink_valid             (mm2stfifo_1_out_valid),                          //       in.valid
		.avalonst_sink_data              (mm2stfifo_1_out_data),                           //         .data
		.avalonst_sink_channel           (mm2stfifo_1_out_channel),                        //         .channel
		.avalonst_sink_error             (mm2stfifo_1_out_error),                          //         .error
		.avalonst_sink_ready             (mm2stfifo_1_out_ready),                          //         .ready
		.avalonmm_read_slave_readdata    (mm_interconnect_0_st2mmfifo_0_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read        (mm_interconnect_0_st2mmfifo_0_out_read),         //         .read
		.avalonmm_read_slave_address     (mm_interconnect_0_st2mmfifo_0_out_address),      //         .address
		.avalonmm_read_slave_waitrequest (mm_interconnect_0_st2mmfifo_0_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address     (mm_interconnect_0_st2mmfifo_0_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read        (mm_interconnect_0_st2mmfifo_0_in_csr_read),      //         .read
		.wrclk_control_slave_writedata   (mm_interconnect_0_st2mmfifo_0_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write       (mm_interconnect_0_st2mmfifo_0_in_csr_write),     //         .write
		.wrclk_control_slave_readdata    (mm_interconnect_0_st2mmfifo_0_in_csr_readdata),  //         .readdata
		.wrclk_control_slave_irq         (irq_mapper_receiver1_irq)                        //   in_irq.irq
	);

	unsaved_ST2MMFIFO_0 st2mmfifo_1 (
		.wrclock                         (clk_clk),                                        //   clk_in.clk
		.reset_n                         (~rst_controller_reset_out_reset),                // reset_in.reset_n
		.avalonst_sink_valid             (mm2stfifo_0_out_valid),                          //       in.valid
		.avalonst_sink_data              (mm2stfifo_0_out_data),                           //         .data
		.avalonst_sink_channel           (mm2stfifo_0_out_channel),                        //         .channel
		.avalonst_sink_error             (mm2stfifo_0_out_error),                          //         .error
		.avalonst_sink_ready             (mm2stfifo_0_out_ready),                          //         .ready
		.avalonmm_read_slave_readdata    (mm_interconnect_0_st2mmfifo_1_out_readdata),     //      out.readdata
		.avalonmm_read_slave_read        (mm_interconnect_0_st2mmfifo_1_out_read),         //         .read
		.avalonmm_read_slave_address     (mm_interconnect_0_st2mmfifo_1_out_address),      //         .address
		.avalonmm_read_slave_waitrequest (mm_interconnect_0_st2mmfifo_1_out_waitrequest),  //         .waitrequest
		.wrclk_control_slave_address     (mm_interconnect_0_st2mmfifo_1_in_csr_address),   //   in_csr.address
		.wrclk_control_slave_read        (mm_interconnect_0_st2mmfifo_1_in_csr_read),      //         .read
		.wrclk_control_slave_writedata   (mm_interconnect_0_st2mmfifo_1_in_csr_writedata), //         .writedata
		.wrclk_control_slave_write       (mm_interconnect_0_st2mmfifo_1_in_csr_write),     //         .write
		.wrclk_control_slave_readdata    (mm_interconnect_0_st2mmfifo_1_in_csr_readdata),  //         .readdata
		.wrclk_control_slave_irq         (irq_mapper_001_receiver1_irq)                    //   in_irq.irq
	);

	unsaved_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver2_irq)                                     //               irq.irq
	);

	unsaved_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (clk_clk),                                                    //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                            //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                         //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                           //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	unsaved_nios2_gen2_1 nios2_gen2_1 (
		.clk                                 (clk_clk),                                                    //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                            //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                         //                          .reset_req
		.d_address                           (nios2_gen2_1_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_1_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_1_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_1_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_1_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_1_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_1_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_1_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_1_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_1_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_1_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_1_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_gen2_1_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                           //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_1_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_1_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_1_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_1_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_1_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_1_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_1_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_1_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	unsaved_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),               //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	unsaved_onchip_memory2_1 onchip_memory2_1 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_1_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_1_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_1_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_1_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_1_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_1_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_1_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),               //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	unsaved_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                  (clk_clk),                                                     //                                clk_0_clk.clk
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                              // nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_data_master_address               (nios2_gen2_0_data_master_address),                            //                 nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest           (nios2_gen2_0_data_master_waitrequest),                        //                                         .waitrequest
		.nios2_gen2_0_data_master_byteenable            (nios2_gen2_0_data_master_byteenable),                         //                                         .byteenable
		.nios2_gen2_0_data_master_read                  (nios2_gen2_0_data_master_read),                               //                                         .read
		.nios2_gen2_0_data_master_readdata              (nios2_gen2_0_data_master_readdata),                           //                                         .readdata
		.nios2_gen2_0_data_master_write                 (nios2_gen2_0_data_master_write),                              //                                         .write
		.nios2_gen2_0_data_master_writedata             (nios2_gen2_0_data_master_writedata),                          //                                         .writedata
		.nios2_gen2_0_data_master_debugaccess           (nios2_gen2_0_data_master_debugaccess),                        //                                         .debugaccess
		.nios2_gen2_0_instruction_master_address        (nios2_gen2_0_instruction_master_address),                     //          nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest    (nios2_gen2_0_instruction_master_waitrequest),                 //                                         .waitrequest
		.nios2_gen2_0_instruction_master_read           (nios2_gen2_0_instruction_master_read),                        //                                         .read
		.nios2_gen2_0_instruction_master_readdata       (nios2_gen2_0_instruction_master_readdata),                    //                                         .readdata
		.nios2_gen2_1_data_master_address               (nios2_gen2_1_data_master_address),                            //                 nios2_gen2_1_data_master.address
		.nios2_gen2_1_data_master_waitrequest           (nios2_gen2_1_data_master_waitrequest),                        //                                         .waitrequest
		.nios2_gen2_1_data_master_byteenable            (nios2_gen2_1_data_master_byteenable),                         //                                         .byteenable
		.nios2_gen2_1_data_master_read                  (nios2_gen2_1_data_master_read),                               //                                         .read
		.nios2_gen2_1_data_master_readdata              (nios2_gen2_1_data_master_readdata),                           //                                         .readdata
		.nios2_gen2_1_data_master_write                 (nios2_gen2_1_data_master_write),                              //                                         .write
		.nios2_gen2_1_data_master_writedata             (nios2_gen2_1_data_master_writedata),                          //                                         .writedata
		.nios2_gen2_1_data_master_debugaccess           (nios2_gen2_1_data_master_debugaccess),                        //                                         .debugaccess
		.nios2_gen2_1_instruction_master_address        (nios2_gen2_1_instruction_master_address),                     //          nios2_gen2_1_instruction_master.address
		.nios2_gen2_1_instruction_master_waitrequest    (nios2_gen2_1_instruction_master_waitrequest),                 //                                         .waitrequest
		.nios2_gen2_1_instruction_master_read           (nios2_gen2_1_instruction_master_read),                        //                                         .read
		.nios2_gen2_1_instruction_master_readdata       (nios2_gen2_1_instruction_master_readdata),                    //                                         .readdata
		.Inst_mem_0_s1_address                          (mm_interconnect_0_inst_mem_0_s1_address),                     //                            Inst_mem_0_s1.address
		.Inst_mem_0_s1_write                            (mm_interconnect_0_inst_mem_0_s1_write),                       //                                         .write
		.Inst_mem_0_s1_readdata                         (mm_interconnect_0_inst_mem_0_s1_readdata),                    //                                         .readdata
		.Inst_mem_0_s1_writedata                        (mm_interconnect_0_inst_mem_0_s1_writedata),                   //                                         .writedata
		.Inst_mem_0_s1_byteenable                       (mm_interconnect_0_inst_mem_0_s1_byteenable),                  //                                         .byteenable
		.Inst_mem_0_s1_chipselect                       (mm_interconnect_0_inst_mem_0_s1_chipselect),                  //                                         .chipselect
		.Inst_mem_0_s1_clken                            (mm_interconnect_0_inst_mem_0_s1_clken),                       //                                         .clken
		.Inst_mem_1_s1_address                          (mm_interconnect_0_inst_mem_1_s1_address),                     //                            Inst_mem_1_s1.address
		.Inst_mem_1_s1_write                            (mm_interconnect_0_inst_mem_1_s1_write),                       //                                         .write
		.Inst_mem_1_s1_readdata                         (mm_interconnect_0_inst_mem_1_s1_readdata),                    //                                         .readdata
		.Inst_mem_1_s1_writedata                        (mm_interconnect_0_inst_mem_1_s1_writedata),                   //                                         .writedata
		.Inst_mem_1_s1_byteenable                       (mm_interconnect_0_inst_mem_1_s1_byteenable),                  //                                         .byteenable
		.Inst_mem_1_s1_chipselect                       (mm_interconnect_0_inst_mem_1_s1_chipselect),                  //                                         .chipselect
		.Inst_mem_1_s1_clken                            (mm_interconnect_0_inst_mem_1_s1_clken),                       //                                         .clken
		.jtag_uart_0_avalon_jtag_slave_address          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //            jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                         .write
		.jtag_uart_0_avalon_jtag_slave_read             (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                         .read
		.jtag_uart_0_avalon_jtag_slave_readdata         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                         .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                         .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest      (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                         .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                         .chipselect
		.MM2STFIFO_0_in_address                         (mm_interconnect_0_mm2stfifo_0_in_address),                    //                           MM2STFIFO_0_in.address
		.MM2STFIFO_0_in_write                           (mm_interconnect_0_mm2stfifo_0_in_write),                      //                                         .write
		.MM2STFIFO_0_in_writedata                       (mm_interconnect_0_mm2stfifo_0_in_writedata),                  //                                         .writedata
		.MM2STFIFO_0_in_waitrequest                     (mm_interconnect_0_mm2stfifo_0_in_waitrequest),                //                                         .waitrequest
		.MM2STFIFO_0_in_csr_address                     (mm_interconnect_0_mm2stfifo_0_in_csr_address),                //                       MM2STFIFO_0_in_csr.address
		.MM2STFIFO_0_in_csr_write                       (mm_interconnect_0_mm2stfifo_0_in_csr_write),                  //                                         .write
		.MM2STFIFO_0_in_csr_read                        (mm_interconnect_0_mm2stfifo_0_in_csr_read),                   //                                         .read
		.MM2STFIFO_0_in_csr_readdata                    (mm_interconnect_0_mm2stfifo_0_in_csr_readdata),               //                                         .readdata
		.MM2STFIFO_0_in_csr_writedata                   (mm_interconnect_0_mm2stfifo_0_in_csr_writedata),              //                                         .writedata
		.MM2STFIFO_1_in_address                         (mm_interconnect_0_mm2stfifo_1_in_address),                    //                           MM2STFIFO_1_in.address
		.MM2STFIFO_1_in_write                           (mm_interconnect_0_mm2stfifo_1_in_write),                      //                                         .write
		.MM2STFIFO_1_in_writedata                       (mm_interconnect_0_mm2stfifo_1_in_writedata),                  //                                         .writedata
		.MM2STFIFO_1_in_waitrequest                     (mm_interconnect_0_mm2stfifo_1_in_waitrequest),                //                                         .waitrequest
		.MM2STFIFO_1_in_csr_address                     (mm_interconnect_0_mm2stfifo_1_in_csr_address),                //                       MM2STFIFO_1_in_csr.address
		.MM2STFIFO_1_in_csr_write                       (mm_interconnect_0_mm2stfifo_1_in_csr_write),                  //                                         .write
		.MM2STFIFO_1_in_csr_read                        (mm_interconnect_0_mm2stfifo_1_in_csr_read),                   //                                         .read
		.MM2STFIFO_1_in_csr_readdata                    (mm_interconnect_0_mm2stfifo_1_in_csr_readdata),               //                                         .readdata
		.MM2STFIFO_1_in_csr_writedata                   (mm_interconnect_0_mm2stfifo_1_in_csr_writedata),              //                                         .writedata
		.nios2_gen2_0_debug_mem_slave_address           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),      //             nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),        //                                         .write
		.nios2_gen2_0_debug_mem_slave_read              (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),         //                                         .read
		.nios2_gen2_0_debug_mem_slave_readdata          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),     //                                         .readdata
		.nios2_gen2_0_debug_mem_slave_writedata         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),    //                                         .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable        (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),   //                                         .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest),  //                                         .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess),  //                                         .debugaccess
		.nios2_gen2_1_debug_mem_slave_address           (mm_interconnect_0_nios2_gen2_1_debug_mem_slave_address),      //             nios2_gen2_1_debug_mem_slave.address
		.nios2_gen2_1_debug_mem_slave_write             (mm_interconnect_0_nios2_gen2_1_debug_mem_slave_write),        //                                         .write
		.nios2_gen2_1_debug_mem_slave_read              (mm_interconnect_0_nios2_gen2_1_debug_mem_slave_read),         //                                         .read
		.nios2_gen2_1_debug_mem_slave_readdata          (mm_interconnect_0_nios2_gen2_1_debug_mem_slave_readdata),     //                                         .readdata
		.nios2_gen2_1_debug_mem_slave_writedata         (mm_interconnect_0_nios2_gen2_1_debug_mem_slave_writedata),    //                                         .writedata
		.nios2_gen2_1_debug_mem_slave_byteenable        (mm_interconnect_0_nios2_gen2_1_debug_mem_slave_byteenable),   //                                         .byteenable
		.nios2_gen2_1_debug_mem_slave_waitrequest       (mm_interconnect_0_nios2_gen2_1_debug_mem_slave_waitrequest),  //                                         .waitrequest
		.nios2_gen2_1_debug_mem_slave_debugaccess       (mm_interconnect_0_nios2_gen2_1_debug_mem_slave_debugaccess),  //                                         .debugaccess
		.onchip_memory2_0_s1_address                    (mm_interconnect_0_onchip_memory2_0_s1_address),               //                      onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                      (mm_interconnect_0_onchip_memory2_0_s1_write),                 //                                         .write
		.onchip_memory2_0_s1_readdata                   (mm_interconnect_0_onchip_memory2_0_s1_readdata),              //                                         .readdata
		.onchip_memory2_0_s1_writedata                  (mm_interconnect_0_onchip_memory2_0_s1_writedata),             //                                         .writedata
		.onchip_memory2_0_s1_byteenable                 (mm_interconnect_0_onchip_memory2_0_s1_byteenable),            //                                         .byteenable
		.onchip_memory2_0_s1_chipselect                 (mm_interconnect_0_onchip_memory2_0_s1_chipselect),            //                                         .chipselect
		.onchip_memory2_0_s1_clken                      (mm_interconnect_0_onchip_memory2_0_s1_clken),                 //                                         .clken
		.onchip_memory2_1_s1_address                    (mm_interconnect_0_onchip_memory2_1_s1_address),               //                      onchip_memory2_1_s1.address
		.onchip_memory2_1_s1_write                      (mm_interconnect_0_onchip_memory2_1_s1_write),                 //                                         .write
		.onchip_memory2_1_s1_readdata                   (mm_interconnect_0_onchip_memory2_1_s1_readdata),              //                                         .readdata
		.onchip_memory2_1_s1_writedata                  (mm_interconnect_0_onchip_memory2_1_s1_writedata),             //                                         .writedata
		.onchip_memory2_1_s1_byteenable                 (mm_interconnect_0_onchip_memory2_1_s1_byteenable),            //                                         .byteenable
		.onchip_memory2_1_s1_chipselect                 (mm_interconnect_0_onchip_memory2_1_s1_chipselect),            //                                         .chipselect
		.onchip_memory2_1_s1_clken                      (mm_interconnect_0_onchip_memory2_1_s1_clken),                 //                                         .clken
		.ST2MMFIFO_0_in_csr_address                     (mm_interconnect_0_st2mmfifo_0_in_csr_address),                //                       ST2MMFIFO_0_in_csr.address
		.ST2MMFIFO_0_in_csr_write                       (mm_interconnect_0_st2mmfifo_0_in_csr_write),                  //                                         .write
		.ST2MMFIFO_0_in_csr_read                        (mm_interconnect_0_st2mmfifo_0_in_csr_read),                   //                                         .read
		.ST2MMFIFO_0_in_csr_readdata                    (mm_interconnect_0_st2mmfifo_0_in_csr_readdata),               //                                         .readdata
		.ST2MMFIFO_0_in_csr_writedata                   (mm_interconnect_0_st2mmfifo_0_in_csr_writedata),              //                                         .writedata
		.ST2MMFIFO_0_out_address                        (mm_interconnect_0_st2mmfifo_0_out_address),                   //                          ST2MMFIFO_0_out.address
		.ST2MMFIFO_0_out_read                           (mm_interconnect_0_st2mmfifo_0_out_read),                      //                                         .read
		.ST2MMFIFO_0_out_readdata                       (mm_interconnect_0_st2mmfifo_0_out_readdata),                  //                                         .readdata
		.ST2MMFIFO_0_out_waitrequest                    (mm_interconnect_0_st2mmfifo_0_out_waitrequest),               //                                         .waitrequest
		.ST2MMFIFO_1_in_csr_address                     (mm_interconnect_0_st2mmfifo_1_in_csr_address),                //                       ST2MMFIFO_1_in_csr.address
		.ST2MMFIFO_1_in_csr_write                       (mm_interconnect_0_st2mmfifo_1_in_csr_write),                  //                                         .write
		.ST2MMFIFO_1_in_csr_read                        (mm_interconnect_0_st2mmfifo_1_in_csr_read),                   //                                         .read
		.ST2MMFIFO_1_in_csr_readdata                    (mm_interconnect_0_st2mmfifo_1_in_csr_readdata),               //                                         .readdata
		.ST2MMFIFO_1_in_csr_writedata                   (mm_interconnect_0_st2mmfifo_1_in_csr_writedata),              //                                         .writedata
		.ST2MMFIFO_1_out_address                        (mm_interconnect_0_st2mmfifo_1_out_address),                   //                          ST2MMFIFO_1_out.address
		.ST2MMFIFO_1_out_read                           (mm_interconnect_0_st2mmfifo_1_out_read),                      //                                         .read
		.ST2MMFIFO_1_out_readdata                       (mm_interconnect_0_st2mmfifo_1_out_readdata),                  //                                         .readdata
		.ST2MMFIFO_1_out_waitrequest                    (mm_interconnect_0_st2mmfifo_1_out_waitrequest)                //                                         .waitrequest
	);

	unsaved_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.sender_irq    (nios2_gen2_0_irq_irq)            //    sender.irq
	);

	unsaved_irq_mapper irq_mapper_001 (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_001_receiver0_irq),   // receiver0.irq
		.receiver1_irq (irq_mapper_001_receiver1_irq),   // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.sender_irq    (nios2_gen2_1_irq_irq)            //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
