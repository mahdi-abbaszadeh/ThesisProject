
module unsaved (
	clk_clk,
	resetn_reset_n);	

	input		clk_clk;
	input		resetn_reset_n;
endmodule
